// Copyright 2024 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Authors:
// - Thomas Benz <tbenz@iis.ee.ethz.ch>
//
// Generated with convert_pcm.py (phsauter@iis.ee.ethz.ch)

module mlem_sound_data #(
    parameter type addr_t = logic
) (
    input  addr_t addr_i,
    output logic  data_o
);
    always_comb begin
        data_o = 1'b0;
        unique case (addr_i)
            0 : data_o = 1'b0;
            1 : data_o = 1'b0;
            2 : data_o = 1'b0;
            3 : data_o = 1'b0;
            4 : data_o = 1'b0;
            5 : data_o = 1'b0;
            6 : data_o = 1'b0;
            7 : data_o = 1'b0;
            8 : data_o = 1'b0;
            9 : data_o = 1'b0;
            10 : data_o = 1'b1;
            11 : data_o = 1'b1;
            12 : data_o = 1'b1;
            13 : data_o = 1'b1;
            14 : data_o = 1'b1;
            15 : data_o = 1'b1;
            16 : data_o = 1'b0;
            17 : data_o = 1'b0;
            18 : data_o = 1'b0;
            19 : data_o = 1'b0;
            20 : data_o = 1'b0;
            21 : data_o = 1'b0;
            22 : data_o = 1'b1;
            23 : data_o = 1'b1;
            24 : data_o = 1'b1;
            25 : data_o = 1'b0;
            26 : data_o = 1'b0;
            27 : data_o = 1'b0;
            28 : data_o = 1'b0;
            29 : data_o = 1'b0;
            30 : data_o = 1'b0;
            31 : data_o = 1'b0;
            32 : data_o = 1'b1;
            33 : data_o = 1'b1;
            34 : data_o = 1'b1;
            35 : data_o = 1'b0;
            36 : data_o = 1'b0;
            37 : data_o = 1'b0;
            38 : data_o = 1'b0;
            39 : data_o = 1'b0;
            40 : data_o = 1'b0;
            41 : data_o = 1'b0;
            42 : data_o = 1'b0;
            43 : data_o = 1'b0;
            44 : data_o = 1'b0;
            45 : data_o = 1'b0;
            46 : data_o = 1'b0;
            47 : data_o = 1'b0;
            48 : data_o = 1'b1;
            49 : data_o = 1'b1;
            50 : data_o = 1'b1;
            51 : data_o = 1'b1;
            52 : data_o = 1'b0;
            53 : data_o = 1'b0;
            54 : data_o = 1'b0;
            55 : data_o = 1'b0;
            56 : data_o = 1'b1;
            57 : data_o = 1'b0;
            58 : data_o = 1'b1;
            59 : data_o = 1'b1;
            60 : data_o = 1'b0;
            61 : data_o = 1'b0;
            62 : data_o = 1'b0;
            63 : data_o = 1'b0;
            64 : data_o = 1'b0;
            65 : data_o = 1'b0;
            66 : data_o = 1'b0;
            67 : data_o = 1'b0;
            68 : data_o = 1'b0;
            69 : data_o = 1'b0;
            70 : data_o = 1'b0;
            71 : data_o = 1'b0;
            72 : data_o = 1'b0;
            73 : data_o = 1'b0;
            74 : data_o = 1'b0;
            75 : data_o = 1'b0;
            76 : data_o = 1'b1;
            77 : data_o = 1'b1;
            78 : data_o = 1'b1;
            79 : data_o = 1'b1;
            80 : data_o = 1'b1;
            81 : data_o = 1'b1;
            82 : data_o = 1'b1;
            83 : data_o = 1'b1;
            84 : data_o = 1'b1;
            85 : data_o = 1'b1;
            86 : data_o = 1'b0;
            87 : data_o = 1'b0;
            88 : data_o = 1'b0;
            89 : data_o = 1'b0;
            90 : data_o = 1'b0;
            91 : data_o = 1'b0;
            92 : data_o = 1'b1;
            93 : data_o = 1'b1;
            94 : data_o = 1'b1;
            95 : data_o = 1'b0;
            96 : data_o = 1'b1;
            97 : data_o = 1'b1;
            98 : data_o = 1'b1;
            99 : data_o = 1'b1;
            100 : data_o = 1'b1;
            101 : data_o = 1'b1;
            102 : data_o = 1'b1;
            103 : data_o = 1'b1;
            104 : data_o = 1'b0;
            105 : data_o = 1'b0;
            106 : data_o = 1'b1;
            107 : data_o = 1'b1;
            108 : data_o = 1'b1;
            109 : data_o = 1'b1;
            110 : data_o = 1'b0;
            111 : data_o = 1'b0;
            112 : data_o = 1'b0;
            113 : data_o = 1'b0;
            114 : data_o = 1'b0;
            115 : data_o = 1'b0;
            116 : data_o = 1'b0;
            117 : data_o = 1'b0;
            118 : data_o = 1'b0;
            119 : data_o = 1'b0;
            120 : data_o = 1'b1;
            121 : data_o = 1'b1;
            122 : data_o = 1'b1;
            123 : data_o = 1'b1;
            124 : data_o = 1'b1;
            125 : data_o = 1'b1;
            126 : data_o = 1'b0;
            127 : data_o = 1'b0;
            128 : data_o = 1'b0;
            129 : data_o = 1'b0;
            130 : data_o = 1'b0;
            131 : data_o = 1'b1;
            132 : data_o = 1'b1;
            133 : data_o = 1'b1;
            134 : data_o = 1'b1;
            135 : data_o = 1'b0;
            136 : data_o = 1'b0;
            137 : data_o = 1'b0;
            138 : data_o = 1'b0;
            139 : data_o = 1'b0;
            140 : data_o = 1'b0;
            141 : data_o = 1'b0;
            142 : data_o = 1'b0;
            143 : data_o = 1'b0;
            144 : data_o = 1'b0;
            145 : data_o = 1'b0;
            146 : data_o = 1'b0;
            147 : data_o = 1'b0;
            148 : data_o = 1'b0;
            149 : data_o = 1'b0;
            150 : data_o = 1'b0;
            151 : data_o = 1'b0;
            152 : data_o = 1'b0;
            153 : data_o = 1'b0;
            154 : data_o = 1'b0;
            155 : data_o = 1'b0;
            156 : data_o = 1'b0;
            157 : data_o = 1'b0;
            158 : data_o = 1'b0;
            159 : data_o = 1'b0;
            160 : data_o = 1'b0;
            161 : data_o = 1'b0;
            162 : data_o = 1'b0;
            163 : data_o = 1'b0;
            164 : data_o = 1'b0;
            165 : data_o = 1'b0;
            166 : data_o = 1'b0;
            167 : data_o = 1'b0;
            168 : data_o = 1'b0;
            169 : data_o = 1'b0;
            170 : data_o = 1'b0;
            171 : data_o = 1'b0;
            172 : data_o = 1'b0;
            173 : data_o = 1'b0;
            174 : data_o = 1'b0;
            175 : data_o = 1'b0;
            176 : data_o = 1'b0;
            177 : data_o = 1'b0;
            178 : data_o = 1'b0;
            179 : data_o = 1'b0;
            180 : data_o = 1'b0;
            181 : data_o = 1'b1;
            182 : data_o = 1'b1;
            183 : data_o = 1'b1;
            184 : data_o = 1'b1;
            185 : data_o = 1'b1;
            186 : data_o = 1'b1;
            187 : data_o = 1'b1;
            188 : data_o = 1'b1;
            189 : data_o = 1'b1;
            190 : data_o = 1'b1;
            191 : data_o = 1'b1;
            192 : data_o = 1'b1;
            193 : data_o = 1'b1;
            194 : data_o = 1'b1;
            195 : data_o = 1'b1;
            196 : data_o = 1'b1;
            197 : data_o = 1'b1;
            198 : data_o = 1'b1;
            199 : data_o = 1'b1;
            200 : data_o = 1'b1;
            201 : data_o = 1'b1;
            202 : data_o = 1'b1;
            203 : data_o = 1'b1;
            204 : data_o = 1'b1;
            205 : data_o = 1'b1;
            206 : data_o = 1'b1;
            207 : data_o = 1'b1;
            208 : data_o = 1'b1;
            209 : data_o = 1'b1;
            210 : data_o = 1'b1;
            211 : data_o = 1'b1;
            212 : data_o = 1'b1;
            213 : data_o = 1'b1;
            214 : data_o = 1'b1;
            215 : data_o = 1'b1;
            216 : data_o = 1'b1;
            217 : data_o = 1'b1;
            218 : data_o = 1'b1;
            219 : data_o = 1'b1;
            220 : data_o = 1'b1;
            221 : data_o = 1'b1;
            222 : data_o = 1'b1;
            223 : data_o = 1'b0;
            224 : data_o = 1'b0;
            225 : data_o = 1'b0;
            226 : data_o = 1'b0;
            227 : data_o = 1'b0;
            228 : data_o = 1'b0;
            229 : data_o = 1'b0;
            230 : data_o = 1'b0;
            231 : data_o = 1'b0;
            232 : data_o = 1'b0;
            233 : data_o = 1'b0;
            234 : data_o = 1'b0;
            235 : data_o = 1'b0;
            236 : data_o = 1'b0;
            237 : data_o = 1'b0;
            238 : data_o = 1'b0;
            239 : data_o = 1'b0;
            240 : data_o = 1'b0;
            241 : data_o = 1'b0;
            242 : data_o = 1'b0;
            243 : data_o = 1'b0;
            244 : data_o = 1'b0;
            245 : data_o = 1'b0;
            246 : data_o = 1'b0;
            247 : data_o = 1'b0;
            248 : data_o = 1'b0;
            249 : data_o = 1'b0;
            250 : data_o = 1'b0;
            251 : data_o = 1'b0;
            252 : data_o = 1'b0;
            253 : data_o = 1'b0;
            254 : data_o = 1'b0;
            255 : data_o = 1'b0;
            256 : data_o = 1'b0;
            257 : data_o = 1'b0;
            258 : data_o = 1'b0;
            259 : data_o = 1'b0;
            260 : data_o = 1'b0;
            261 : data_o = 1'b0;
            262 : data_o = 1'b1;
            263 : data_o = 1'b1;
            264 : data_o = 1'b1;
            265 : data_o = 1'b1;
            266 : data_o = 1'b1;
            267 : data_o = 1'b1;
            268 : data_o = 1'b1;
            269 : data_o = 1'b1;
            270 : data_o = 1'b1;
            271 : data_o = 1'b1;
            272 : data_o = 1'b1;
            273 : data_o = 1'b1;
            274 : data_o = 1'b1;
            275 : data_o = 1'b0;
            276 : data_o = 1'b0;
            277 : data_o = 1'b0;
            278 : data_o = 1'b0;
            279 : data_o = 1'b0;
            280 : data_o = 1'b0;
            281 : data_o = 1'b0;
            282 : data_o = 1'b0;
            283 : data_o = 1'b0;
            284 : data_o = 1'b0;
            285 : data_o = 1'b0;
            286 : data_o = 1'b0;
            287 : data_o = 1'b0;
            288 : data_o = 1'b0;
            289 : data_o = 1'b0;
            290 : data_o = 1'b0;
            291 : data_o = 1'b0;
            292 : data_o = 1'b0;
            293 : data_o = 1'b1;
            294 : data_o = 1'b1;
            295 : data_o = 1'b1;
            296 : data_o = 1'b1;
            297 : data_o = 1'b1;
            298 : data_o = 1'b1;
            299 : data_o = 1'b1;
            300 : data_o = 1'b1;
            301 : data_o = 1'b1;
            302 : data_o = 1'b1;
            303 : data_o = 1'b1;
            304 : data_o = 1'b1;
            305 : data_o = 1'b1;
            306 : data_o = 1'b1;
            307 : data_o = 1'b1;
            308 : data_o = 1'b1;
            309 : data_o = 1'b1;
            310 : data_o = 1'b1;
            311 : data_o = 1'b1;
            312 : data_o = 1'b1;
            313 : data_o = 1'b1;
            314 : data_o = 1'b1;
            315 : data_o = 1'b1;
            316 : data_o = 1'b1;
            317 : data_o = 1'b1;
            318 : data_o = 1'b1;
            319 : data_o = 1'b1;
            320 : data_o = 1'b1;
            321 : data_o = 1'b1;
            322 : data_o = 1'b1;
            323 : data_o = 1'b1;
            324 : data_o = 1'b0;
            325 : data_o = 1'b0;
            326 : data_o = 1'b0;
            327 : data_o = 1'b0;
            328 : data_o = 1'b0;
            329 : data_o = 1'b1;
            330 : data_o = 1'b1;
            331 : data_o = 1'b1;
            332 : data_o = 1'b1;
            333 : data_o = 1'b0;
            334 : data_o = 1'b0;
            335 : data_o = 1'b0;
            336 : data_o = 1'b0;
            337 : data_o = 1'b0;
            338 : data_o = 1'b0;
            339 : data_o = 1'b0;
            340 : data_o = 1'b0;
            341 : data_o = 1'b0;
            342 : data_o = 1'b0;
            343 : data_o = 1'b0;
            344 : data_o = 1'b0;
            345 : data_o = 1'b0;
            346 : data_o = 1'b0;
            347 : data_o = 1'b0;
            348 : data_o = 1'b0;
            349 : data_o = 1'b0;
            350 : data_o = 1'b0;
            351 : data_o = 1'b0;
            352 : data_o = 1'b0;
            353 : data_o = 1'b0;
            354 : data_o = 1'b0;
            355 : data_o = 1'b0;
            356 : data_o = 1'b0;
            357 : data_o = 1'b0;
            358 : data_o = 1'b0;
            359 : data_o = 1'b0;
            360 : data_o = 1'b0;
            361 : data_o = 1'b0;
            362 : data_o = 1'b1;
            363 : data_o = 1'b1;
            364 : data_o = 1'b1;
            365 : data_o = 1'b1;
            366 : data_o = 1'b1;
            367 : data_o = 1'b0;
            368 : data_o = 1'b0;
            369 : data_o = 1'b0;
            370 : data_o = 1'b0;
            371 : data_o = 1'b0;
            372 : data_o = 1'b1;
            373 : data_o = 1'b1;
            374 : data_o = 1'b1;
            375 : data_o = 1'b1;
            376 : data_o = 1'b1;
            377 : data_o = 1'b1;
            378 : data_o = 1'b1;
            379 : data_o = 1'b1;
            380 : data_o = 1'b1;
            381 : data_o = 1'b1;
            382 : data_o = 1'b1;
            383 : data_o = 1'b1;
            384 : data_o = 1'b1;
            385 : data_o = 1'b1;
            386 : data_o = 1'b1;
            387 : data_o = 1'b1;
            388 : data_o = 1'b1;
            389 : data_o = 1'b1;
            390 : data_o = 1'b1;
            391 : data_o = 1'b1;
            392 : data_o = 1'b1;
            393 : data_o = 1'b1;
            394 : data_o = 1'b1;
            395 : data_o = 1'b1;
            396 : data_o = 1'b1;
            397 : data_o = 1'b1;
            398 : data_o = 1'b1;
            399 : data_o = 1'b1;
            400 : data_o = 1'b0;
            401 : data_o = 1'b0;
            402 : data_o = 1'b0;
            403 : data_o = 1'b0;
            404 : data_o = 1'b0;
            405 : data_o = 1'b0;
            406 : data_o = 1'b0;
            407 : data_o = 1'b0;
            408 : data_o = 1'b0;
            409 : data_o = 1'b0;
            410 : data_o = 1'b0;
            411 : data_o = 1'b1;
            412 : data_o = 1'b1;
            413 : data_o = 1'b1;
            414 : data_o = 1'b1;
            415 : data_o = 1'b1;
            416 : data_o = 1'b1;
            417 : data_o = 1'b1;
            418 : data_o = 1'b1;
            419 : data_o = 1'b1;
            420 : data_o = 1'b1;
            421 : data_o = 1'b1;
            422 : data_o = 1'b1;
            423 : data_o = 1'b1;
            424 : data_o = 1'b1;
            425 : data_o = 1'b1;
            426 : data_o = 1'b1;
            427 : data_o = 1'b1;
            428 : data_o = 1'b1;
            429 : data_o = 1'b1;
            430 : data_o = 1'b1;
            431 : data_o = 1'b1;
            432 : data_o = 1'b1;
            433 : data_o = 1'b0;
            434 : data_o = 1'b0;
            435 : data_o = 1'b0;
            436 : data_o = 1'b0;
            437 : data_o = 1'b0;
            438 : data_o = 1'b0;
            439 : data_o = 1'b0;
            440 : data_o = 1'b0;
            441 : data_o = 1'b0;
            442 : data_o = 1'b0;
            443 : data_o = 1'b0;
            444 : data_o = 1'b0;
            445 : data_o = 1'b0;
            446 : data_o = 1'b0;
            447 : data_o = 1'b0;
            448 : data_o = 1'b0;
            449 : data_o = 1'b0;
            450 : data_o = 1'b0;
            451 : data_o = 1'b0;
            452 : data_o = 1'b0;
            453 : data_o = 1'b0;
            454 : data_o = 1'b0;
            455 : data_o = 1'b0;
            456 : data_o = 1'b0;
            457 : data_o = 1'b0;
            458 : data_o = 1'b0;
            459 : data_o = 1'b0;
            460 : data_o = 1'b0;
            461 : data_o = 1'b0;
            462 : data_o = 1'b0;
            463 : data_o = 1'b0;
            464 : data_o = 1'b0;
            465 : data_o = 1'b0;
            466 : data_o = 1'b0;
            467 : data_o = 1'b0;
            468 : data_o = 1'b0;
            469 : data_o = 1'b0;
            470 : data_o = 1'b0;
            471 : data_o = 1'b0;
            472 : data_o = 1'b0;
            473 : data_o = 1'b0;
            474 : data_o = 1'b0;
            475 : data_o = 1'b0;
            476 : data_o = 1'b0;
            477 : data_o = 1'b0;
            478 : data_o = 1'b0;
            479 : data_o = 1'b0;
            480 : data_o = 1'b0;
            481 : data_o = 1'b0;
            482 : data_o = 1'b1;
            483 : data_o = 1'b1;
            484 : data_o = 1'b1;
            485 : data_o = 1'b1;
            486 : data_o = 1'b0;
            487 : data_o = 1'b0;
            488 : data_o = 1'b0;
            489 : data_o = 1'b0;
            490 : data_o = 1'b0;
            491 : data_o = 1'b0;
            492 : data_o = 1'b0;
            493 : data_o = 1'b0;
            494 : data_o = 1'b0;
            495 : data_o = 1'b0;
            496 : data_o = 1'b0;
            497 : data_o = 1'b0;
            498 : data_o = 1'b0;
            499 : data_o = 1'b1;
            500 : data_o = 1'b1;
            501 : data_o = 1'b1;
            502 : data_o = 1'b1;
            503 : data_o = 1'b1;
            504 : data_o = 1'b1;
            505 : data_o = 1'b1;
            506 : data_o = 1'b1;
            507 : data_o = 1'b1;
            508 : data_o = 1'b1;
            509 : data_o = 1'b1;
            510 : data_o = 1'b1;
            511 : data_o = 1'b1;
            512 : data_o = 1'b1;
            513 : data_o = 1'b1;
            514 : data_o = 1'b1;
            515 : data_o = 1'b1;
            516 : data_o = 1'b1;
            517 : data_o = 1'b1;
            518 : data_o = 1'b1;
            519 : data_o = 1'b1;
            520 : data_o = 1'b1;
            521 : data_o = 1'b1;
            522 : data_o = 1'b1;
            523 : data_o = 1'b0;
            524 : data_o = 1'b0;
            525 : data_o = 1'b0;
            526 : data_o = 1'b0;
            527 : data_o = 1'b0;
            528 : data_o = 1'b0;
            529 : data_o = 1'b0;
            530 : data_o = 1'b0;
            531 : data_o = 1'b0;
            532 : data_o = 1'b0;
            533 : data_o = 1'b0;
            534 : data_o = 1'b1;
            535 : data_o = 1'b1;
            536 : data_o = 1'b1;
            537 : data_o = 1'b1;
            538 : data_o = 1'b1;
            539 : data_o = 1'b1;
            540 : data_o = 1'b1;
            541 : data_o = 1'b1;
            542 : data_o = 1'b1;
            543 : data_o = 1'b1;
            544 : data_o = 1'b1;
            545 : data_o = 1'b1;
            546 : data_o = 1'b1;
            547 : data_o = 1'b1;
            548 : data_o = 1'b1;
            549 : data_o = 1'b1;
            550 : data_o = 1'b1;
            551 : data_o = 1'b1;
            552 : data_o = 1'b1;
            553 : data_o = 1'b0;
            554 : data_o = 1'b0;
            555 : data_o = 1'b0;
            556 : data_o = 1'b0;
            557 : data_o = 1'b0;
            558 : data_o = 1'b0;
            559 : data_o = 1'b0;
            560 : data_o = 1'b0;
            561 : data_o = 1'b0;
            562 : data_o = 1'b0;
            563 : data_o = 1'b0;
            564 : data_o = 1'b0;
            565 : data_o = 1'b0;
            566 : data_o = 1'b0;
            567 : data_o = 1'b0;
            568 : data_o = 1'b0;
            569 : data_o = 1'b0;
            570 : data_o = 1'b0;
            571 : data_o = 1'b0;
            572 : data_o = 1'b1;
            573 : data_o = 1'b1;
            574 : data_o = 1'b1;
            575 : data_o = 1'b1;
            576 : data_o = 1'b1;
            577 : data_o = 1'b1;
            578 : data_o = 1'b1;
            579 : data_o = 1'b1;
            580 : data_o = 1'b1;
            581 : data_o = 1'b1;
            582 : data_o = 1'b1;
            583 : data_o = 1'b1;
            584 : data_o = 1'b1;
            585 : data_o = 1'b0;
            586 : data_o = 1'b0;
            587 : data_o = 1'b0;
            588 : data_o = 1'b0;
            589 : data_o = 1'b0;
            590 : data_o = 1'b0;
            591 : data_o = 1'b0;
            592 : data_o = 1'b0;
            593 : data_o = 1'b0;
            594 : data_o = 1'b0;
            595 : data_o = 1'b0;
            596 : data_o = 1'b0;
            597 : data_o = 1'b0;
            598 : data_o = 1'b0;
            599 : data_o = 1'b0;
            600 : data_o = 1'b0;
            601 : data_o = 1'b0;
            602 : data_o = 1'b0;
            603 : data_o = 1'b0;
            604 : data_o = 1'b0;
            605 : data_o = 1'b0;
            606 : data_o = 1'b0;
            607 : data_o = 1'b0;
            608 : data_o = 1'b0;
            609 : data_o = 1'b0;
            610 : data_o = 1'b0;
            611 : data_o = 1'b0;
            612 : data_o = 1'b0;
            613 : data_o = 1'b0;
            614 : data_o = 1'b0;
            615 : data_o = 1'b0;
            616 : data_o = 1'b0;
            617 : data_o = 1'b0;
            618 : data_o = 1'b0;
            619 : data_o = 1'b0;
            620 : data_o = 1'b0;
            621 : data_o = 1'b0;
            622 : data_o = 1'b0;
            623 : data_o = 1'b0;
            624 : data_o = 1'b0;
            625 : data_o = 1'b0;
            626 : data_o = 1'b1;
            627 : data_o = 1'b1;
            628 : data_o = 1'b1;
            629 : data_o = 1'b1;
            630 : data_o = 1'b1;
            631 : data_o = 1'b1;
            632 : data_o = 1'b1;
            633 : data_o = 1'b1;
            634 : data_o = 1'b1;
            635 : data_o = 1'b1;
            636 : data_o = 1'b1;
            637 : data_o = 1'b1;
            638 : data_o = 1'b1;
            639 : data_o = 1'b1;
            640 : data_o = 1'b1;
            641 : data_o = 1'b1;
            642 : data_o = 1'b1;
            643 : data_o = 1'b1;
            644 : data_o = 1'b1;
            645 : data_o = 1'b1;
            646 : data_o = 1'b1;
            647 : data_o = 1'b0;
            648 : data_o = 1'b0;
            649 : data_o = 1'b0;
            650 : data_o = 1'b0;
            651 : data_o = 1'b0;
            652 : data_o = 1'b0;
            653 : data_o = 1'b0;
            654 : data_o = 1'b0;
            655 : data_o = 1'b0;
            656 : data_o = 1'b0;
            657 : data_o = 1'b0;
            658 : data_o = 1'b0;
            659 : data_o = 1'b0;
            660 : data_o = 1'b0;
            661 : data_o = 1'b1;
            662 : data_o = 1'b1;
            663 : data_o = 1'b1;
            664 : data_o = 1'b1;
            665 : data_o = 1'b1;
            666 : data_o = 1'b1;
            667 : data_o = 1'b1;
            668 : data_o = 1'b1;
            669 : data_o = 1'b1;
            670 : data_o = 1'b1;
            671 : data_o = 1'b1;
            672 : data_o = 1'b1;
            673 : data_o = 1'b1;
            674 : data_o = 1'b1;
            675 : data_o = 1'b1;
            676 : data_o = 1'b1;
            677 : data_o = 1'b1;
            678 : data_o = 1'b0;
            679 : data_o = 1'b0;
            680 : data_o = 1'b0;
            681 : data_o = 1'b0;
            682 : data_o = 1'b0;
            683 : data_o = 1'b0;
            684 : data_o = 1'b0;
            685 : data_o = 1'b0;
            686 : data_o = 1'b0;
            687 : data_o = 1'b0;
            688 : data_o = 1'b0;
            689 : data_o = 1'b0;
            690 : data_o = 1'b0;
            691 : data_o = 1'b1;
            692 : data_o = 1'b1;
            693 : data_o = 1'b1;
            694 : data_o = 1'b1;
            695 : data_o = 1'b1;
            696 : data_o = 1'b1;
            697 : data_o = 1'b1;
            698 : data_o = 1'b1;
            699 : data_o = 1'b1;
            700 : data_o = 1'b1;
            701 : data_o = 1'b1;
            702 : data_o = 1'b1;
            703 : data_o = 1'b1;
            704 : data_o = 1'b1;
            705 : data_o = 1'b1;
            706 : data_o = 1'b1;
            707 : data_o = 1'b1;
            708 : data_o = 1'b1;
            709 : data_o = 1'b1;
            710 : data_o = 1'b0;
            711 : data_o = 1'b0;
            712 : data_o = 1'b0;
            713 : data_o = 1'b0;
            714 : data_o = 1'b0;
            715 : data_o = 1'b0;
            716 : data_o = 1'b0;
            717 : data_o = 1'b0;
            718 : data_o = 1'b0;
            719 : data_o = 1'b0;
            720 : data_o = 1'b0;
            721 : data_o = 1'b0;
            722 : data_o = 1'b0;
            723 : data_o = 1'b0;
            724 : data_o = 1'b0;
            725 : data_o = 1'b0;
            726 : data_o = 1'b0;
            727 : data_o = 1'b0;
            728 : data_o = 1'b0;
            729 : data_o = 1'b0;
            730 : data_o = 1'b0;
            731 : data_o = 1'b0;
            732 : data_o = 1'b0;
            733 : data_o = 1'b0;
            734 : data_o = 1'b0;
            735 : data_o = 1'b0;
            736 : data_o = 1'b0;
            737 : data_o = 1'b0;
            738 : data_o = 1'b0;
            739 : data_o = 1'b0;
            740 : data_o = 1'b0;
            741 : data_o = 1'b0;
            742 : data_o = 1'b0;
            743 : data_o = 1'b0;
            744 : data_o = 1'b0;
            745 : data_o = 1'b0;
            746 : data_o = 1'b0;
            747 : data_o = 1'b0;
            748 : data_o = 1'b0;
            749 : data_o = 1'b0;
            750 : data_o = 1'b0;
            751 : data_o = 1'b0;
            752 : data_o = 1'b0;
            753 : data_o = 1'b1;
            754 : data_o = 1'b1;
            755 : data_o = 1'b1;
            756 : data_o = 1'b1;
            757 : data_o = 1'b1;
            758 : data_o = 1'b1;
            759 : data_o = 1'b1;
            760 : data_o = 1'b1;
            761 : data_o = 1'b1;
            762 : data_o = 1'b1;
            763 : data_o = 1'b1;
            764 : data_o = 1'b1;
            765 : data_o = 1'b1;
            766 : data_o = 1'b1;
            767 : data_o = 1'b1;
            768 : data_o = 1'b1;
            769 : data_o = 1'b1;
            770 : data_o = 1'b1;
            771 : data_o = 1'b1;
            772 : data_o = 1'b1;
            773 : data_o = 1'b0;
            774 : data_o = 1'b0;
            775 : data_o = 1'b0;
            776 : data_o = 1'b0;
            777 : data_o = 1'b0;
            778 : data_o = 1'b0;
            779 : data_o = 1'b0;
            780 : data_o = 1'b0;
            781 : data_o = 1'b0;
            782 : data_o = 1'b0;
            783 : data_o = 1'b0;
            784 : data_o = 1'b0;
            785 : data_o = 1'b0;
            786 : data_o = 1'b0;
            787 : data_o = 1'b1;
            788 : data_o = 1'b1;
            789 : data_o = 1'b1;
            790 : data_o = 1'b1;
            791 : data_o = 1'b1;
            792 : data_o = 1'b1;
            793 : data_o = 1'b1;
            794 : data_o = 1'b1;
            795 : data_o = 1'b1;
            796 : data_o = 1'b1;
            797 : data_o = 1'b1;
            798 : data_o = 1'b1;
            799 : data_o = 1'b1;
            800 : data_o = 1'b1;
            801 : data_o = 1'b1;
            802 : data_o = 1'b0;
            803 : data_o = 1'b0;
            804 : data_o = 1'b0;
            805 : data_o = 1'b0;
            806 : data_o = 1'b0;
            807 : data_o = 1'b0;
            808 : data_o = 1'b0;
            809 : data_o = 1'b0;
            810 : data_o = 1'b0;
            811 : data_o = 1'b0;
            812 : data_o = 1'b0;
            813 : data_o = 1'b0;
            814 : data_o = 1'b0;
            815 : data_o = 1'b0;
            816 : data_o = 1'b1;
            817 : data_o = 1'b1;
            818 : data_o = 1'b1;
            819 : data_o = 1'b1;
            820 : data_o = 1'b1;
            821 : data_o = 1'b1;
            822 : data_o = 1'b1;
            823 : data_o = 1'b1;
            824 : data_o = 1'b1;
            825 : data_o = 1'b1;
            826 : data_o = 1'b1;
            827 : data_o = 1'b1;
            828 : data_o = 1'b1;
            829 : data_o = 1'b1;
            830 : data_o = 1'b1;
            831 : data_o = 1'b1;
            832 : data_o = 1'b1;
            833 : data_o = 1'b1;
            834 : data_o = 1'b1;
            835 : data_o = 1'b1;
            836 : data_o = 1'b1;
            837 : data_o = 1'b0;
            838 : data_o = 1'b0;
            839 : data_o = 1'b0;
            840 : data_o = 1'b0;
            841 : data_o = 1'b0;
            842 : data_o = 1'b0;
            843 : data_o = 1'b0;
            844 : data_o = 1'b0;
            845 : data_o = 1'b0;
            846 : data_o = 1'b0;
            847 : data_o = 1'b0;
            848 : data_o = 1'b0;
            849 : data_o = 1'b0;
            850 : data_o = 1'b0;
            851 : data_o = 1'b0;
            852 : data_o = 1'b0;
            853 : data_o = 1'b0;
            854 : data_o = 1'b0;
            855 : data_o = 1'b0;
            856 : data_o = 1'b0;
            857 : data_o = 1'b0;
            858 : data_o = 1'b0;
            859 : data_o = 1'b0;
            860 : data_o = 1'b0;
            861 : data_o = 1'b0;
            862 : data_o = 1'b0;
            863 : data_o = 1'b0;
            864 : data_o = 1'b0;
            865 : data_o = 1'b0;
            866 : data_o = 1'b0;
            867 : data_o = 1'b0;
            868 : data_o = 1'b0;
            869 : data_o = 1'b0;
            870 : data_o = 1'b0;
            871 : data_o = 1'b0;
            872 : data_o = 1'b0;
            873 : data_o = 1'b0;
            874 : data_o = 1'b0;
            875 : data_o = 1'b0;
            876 : data_o = 1'b0;
            877 : data_o = 1'b0;
            878 : data_o = 1'b1;
            879 : data_o = 1'b1;
            880 : data_o = 1'b1;
            881 : data_o = 1'b1;
            882 : data_o = 1'b1;
            883 : data_o = 1'b1;
            884 : data_o = 1'b1;
            885 : data_o = 1'b1;
            886 : data_o = 1'b1;
            887 : data_o = 1'b1;
            888 : data_o = 1'b1;
            889 : data_o = 1'b1;
            890 : data_o = 1'b1;
            891 : data_o = 1'b1;
            892 : data_o = 1'b1;
            893 : data_o = 1'b1;
            894 : data_o = 1'b1;
            895 : data_o = 1'b1;
            896 : data_o = 1'b1;
            897 : data_o = 1'b1;
            898 : data_o = 1'b0;
            899 : data_o = 1'b0;
            900 : data_o = 1'b0;
            901 : data_o = 1'b0;
            902 : data_o = 1'b0;
            903 : data_o = 1'b0;
            904 : data_o = 1'b0;
            905 : data_o = 1'b0;
            906 : data_o = 1'b0;
            907 : data_o = 1'b0;
            908 : data_o = 1'b1;
            909 : data_o = 1'b1;
            910 : data_o = 1'b1;
            911 : data_o = 1'b1;
            912 : data_o = 1'b1;
            913 : data_o = 1'b1;
            914 : data_o = 1'b1;
            915 : data_o = 1'b1;
            916 : data_o = 1'b1;
            917 : data_o = 1'b1;
            918 : data_o = 1'b1;
            919 : data_o = 1'b1;
            920 : data_o = 1'b1;
            921 : data_o = 1'b1;
            922 : data_o = 1'b1;
            923 : data_o = 1'b1;
            924 : data_o = 1'b1;
            925 : data_o = 1'b1;
            926 : data_o = 1'b0;
            927 : data_o = 1'b0;
            928 : data_o = 1'b0;
            929 : data_o = 1'b0;
            930 : data_o = 1'b0;
            931 : data_o = 1'b0;
            932 : data_o = 1'b0;
            933 : data_o = 1'b0;
            934 : data_o = 1'b0;
            935 : data_o = 1'b0;
            936 : data_o = 1'b0;
            937 : data_o = 1'b0;
            938 : data_o = 1'b0;
            939 : data_o = 1'b0;
            940 : data_o = 1'b0;
            941 : data_o = 1'b1;
            942 : data_o = 1'b1;
            943 : data_o = 1'b1;
            944 : data_o = 1'b1;
            945 : data_o = 1'b1;
            946 : data_o = 1'b1;
            947 : data_o = 1'b1;
            948 : data_o = 1'b1;
            949 : data_o = 1'b1;
            950 : data_o = 1'b1;
            951 : data_o = 1'b1;
            952 : data_o = 1'b1;
            953 : data_o = 1'b1;
            954 : data_o = 1'b1;
            955 : data_o = 1'b1;
            956 : data_o = 1'b1;
            957 : data_o = 1'b1;
            958 : data_o = 1'b1;
            959 : data_o = 1'b1;
            960 : data_o = 1'b1;
            961 : data_o = 1'b1;
            962 : data_o = 1'b1;
            963 : data_o = 1'b1;
            964 : data_o = 1'b0;
            965 : data_o = 1'b0;
            966 : data_o = 1'b0;
            967 : data_o = 1'b0;
            968 : data_o = 1'b0;
            969 : data_o = 1'b0;
            970 : data_o = 1'b0;
            971 : data_o = 1'b0;
            972 : data_o = 1'b0;
            973 : data_o = 1'b0;
            974 : data_o = 1'b0;
            975 : data_o = 1'b0;
            976 : data_o = 1'b0;
            977 : data_o = 1'b0;
            978 : data_o = 1'b0;
            979 : data_o = 1'b0;
            980 : data_o = 1'b1;
            981 : data_o = 1'b0;
            982 : data_o = 1'b0;
            983 : data_o = 1'b0;
            984 : data_o = 1'b0;
            985 : data_o = 1'b0;
            986 : data_o = 1'b0;
            987 : data_o = 1'b0;
            988 : data_o = 1'b0;
            989 : data_o = 1'b0;
            990 : data_o = 1'b0;
            991 : data_o = 1'b0;
            992 : data_o = 1'b0;
            993 : data_o = 1'b0;
            994 : data_o = 1'b0;
            995 : data_o = 1'b0;
            996 : data_o = 1'b0;
            997 : data_o = 1'b0;
            998 : data_o = 1'b0;
            999 : data_o = 1'b0;
            1000 : data_o = 1'b0;
            1001 : data_o = 1'b0;
            1002 : data_o = 1'b0;
            1003 : data_o = 1'b1;
            1004 : data_o = 1'b1;
            1005 : data_o = 1'b1;
            1006 : data_o = 1'b1;
            1007 : data_o = 1'b1;
            1008 : data_o = 1'b1;
            1009 : data_o = 1'b1;
            1010 : data_o = 1'b1;
            1011 : data_o = 1'b1;
            1012 : data_o = 1'b1;
            1013 : data_o = 1'b1;
            1014 : data_o = 1'b1;
            1015 : data_o = 1'b1;
            1016 : data_o = 1'b1;
            1017 : data_o = 1'b1;
            1018 : data_o = 1'b0;
            1019 : data_o = 1'b0;
            1020 : data_o = 1'b0;
            1021 : data_o = 1'b0;
            1022 : data_o = 1'b0;
            1023 : data_o = 1'b0;
            1024 : data_o = 1'b0;
            1025 : data_o = 1'b0;
            1026 : data_o = 1'b0;
            1027 : data_o = 1'b0;
            1028 : data_o = 1'b0;
            1029 : data_o = 1'b0;
            1030 : data_o = 1'b0;
            1031 : data_o = 1'b0;
            1032 : data_o = 1'b1;
            1033 : data_o = 1'b1;
            1034 : data_o = 1'b1;
            1035 : data_o = 1'b1;
            1036 : data_o = 1'b1;
            1037 : data_o = 1'b1;
            1038 : data_o = 1'b1;
            1039 : data_o = 1'b1;
            1040 : data_o = 1'b1;
            1041 : data_o = 1'b1;
            1042 : data_o = 1'b1;
            1043 : data_o = 1'b1;
            1044 : data_o = 1'b1;
            1045 : data_o = 1'b1;
            1046 : data_o = 1'b1;
            1047 : data_o = 1'b0;
            1048 : data_o = 1'b0;
            1049 : data_o = 1'b0;
            1050 : data_o = 1'b0;
            1051 : data_o = 1'b0;
            1052 : data_o = 1'b0;
            1053 : data_o = 1'b0;
            1054 : data_o = 1'b0;
            1055 : data_o = 1'b0;
            1056 : data_o = 1'b0;
            1057 : data_o = 1'b0;
            1058 : data_o = 1'b0;
            1059 : data_o = 1'b0;
            1060 : data_o = 1'b0;
            1061 : data_o = 1'b1;
            1062 : data_o = 1'b1;
            1063 : data_o = 1'b1;
            1064 : data_o = 1'b1;
            1065 : data_o = 1'b1;
            1066 : data_o = 1'b1;
            1067 : data_o = 1'b1;
            1068 : data_o = 1'b1;
            1069 : data_o = 1'b1;
            1070 : data_o = 1'b1;
            1071 : data_o = 1'b1;
            1072 : data_o = 1'b1;
            1073 : data_o = 1'b1;
            1074 : data_o = 1'b1;
            1075 : data_o = 1'b1;
            1076 : data_o = 1'b1;
            1077 : data_o = 1'b0;
            1078 : data_o = 1'b1;
            1079 : data_o = 1'b1;
            1080 : data_o = 1'b1;
            1081 : data_o = 1'b1;
            1082 : data_o = 1'b1;
            1083 : data_o = 1'b0;
            1084 : data_o = 1'b0;
            1085 : data_o = 1'b0;
            1086 : data_o = 1'b0;
            1087 : data_o = 1'b0;
            1088 : data_o = 1'b0;
            1089 : data_o = 1'b0;
            1090 : data_o = 1'b0;
            1091 : data_o = 1'b0;
            1092 : data_o = 1'b0;
            1093 : data_o = 1'b0;
            1094 : data_o = 1'b0;
            1095 : data_o = 1'b0;
            1096 : data_o = 1'b0;
            1097 : data_o = 1'b0;
            1098 : data_o = 1'b0;
            1099 : data_o = 1'b0;
            1100 : data_o = 1'b0;
            1101 : data_o = 1'b0;
            1102 : data_o = 1'b0;
            1103 : data_o = 1'b0;
            1104 : data_o = 1'b0;
            1105 : data_o = 1'b0;
            1106 : data_o = 1'b0;
            1107 : data_o = 1'b0;
            1108 : data_o = 1'b0;
            1109 : data_o = 1'b0;
            1110 : data_o = 1'b0;
            1111 : data_o = 1'b0;
            1112 : data_o = 1'b0;
            1113 : data_o = 1'b0;
            1114 : data_o = 1'b0;
            1115 : data_o = 1'b0;
            1116 : data_o = 1'b0;
            1117 : data_o = 1'b0;
            1118 : data_o = 1'b0;
            1119 : data_o = 1'b0;
            1120 : data_o = 1'b0;
            1121 : data_o = 1'b0;
            1122 : data_o = 1'b0;
            1123 : data_o = 1'b0;
            1124 : data_o = 1'b0;
            1125 : data_o = 1'b0;
            1126 : data_o = 1'b0;
            1127 : data_o = 1'b0;
            1128 : data_o = 1'b1;
            1129 : data_o = 1'b1;
            1130 : data_o = 1'b1;
            1131 : data_o = 1'b1;
            1132 : data_o = 1'b1;
            1133 : data_o = 1'b1;
            1134 : data_o = 1'b1;
            1135 : data_o = 1'b1;
            1136 : data_o = 1'b1;
            1137 : data_o = 1'b1;
            1138 : data_o = 1'b1;
            1139 : data_o = 1'b1;
            1140 : data_o = 1'b1;
            1141 : data_o = 1'b1;
            1142 : data_o = 1'b1;
            1143 : data_o = 1'b1;
            1144 : data_o = 1'b0;
            1145 : data_o = 1'b0;
            1146 : data_o = 1'b0;
            1147 : data_o = 1'b0;
            1148 : data_o = 1'b0;
            1149 : data_o = 1'b0;
            1150 : data_o = 1'b0;
            1151 : data_o = 1'b0;
            1152 : data_o = 1'b0;
            1153 : data_o = 1'b0;
            1154 : data_o = 1'b0;
            1155 : data_o = 1'b0;
            1156 : data_o = 1'b0;
            1157 : data_o = 1'b1;
            1158 : data_o = 1'b1;
            1159 : data_o = 1'b1;
            1160 : data_o = 1'b1;
            1161 : data_o = 1'b1;
            1162 : data_o = 1'b1;
            1163 : data_o = 1'b1;
            1164 : data_o = 1'b1;
            1165 : data_o = 1'b1;
            1166 : data_o = 1'b1;
            1167 : data_o = 1'b1;
            1168 : data_o = 1'b1;
            1169 : data_o = 1'b1;
            1170 : data_o = 1'b1;
            1171 : data_o = 1'b1;
            1172 : data_o = 1'b1;
            1173 : data_o = 1'b0;
            1174 : data_o = 1'b0;
            1175 : data_o = 1'b0;
            1176 : data_o = 1'b0;
            1177 : data_o = 1'b0;
            1178 : data_o = 1'b0;
            1179 : data_o = 1'b0;
            1180 : data_o = 1'b0;
            1181 : data_o = 1'b0;
            1182 : data_o = 1'b0;
            1183 : data_o = 1'b0;
            1184 : data_o = 1'b0;
            1185 : data_o = 1'b0;
            1186 : data_o = 1'b1;
            1187 : data_o = 1'b1;
            1188 : data_o = 1'b1;
            1189 : data_o = 1'b1;
            1190 : data_o = 1'b1;
            1191 : data_o = 1'b1;
            1192 : data_o = 1'b1;
            1193 : data_o = 1'b1;
            1194 : data_o = 1'b1;
            1195 : data_o = 1'b1;
            1196 : data_o = 1'b1;
            1197 : data_o = 1'b1;
            1198 : data_o = 1'b1;
            1199 : data_o = 1'b1;
            1200 : data_o = 1'b1;
            1201 : data_o = 1'b0;
            1202 : data_o = 1'b0;
            1203 : data_o = 1'b0;
            1204 : data_o = 1'b0;
            1205 : data_o = 1'b0;
            1206 : data_o = 1'b1;
            1207 : data_o = 1'b1;
            1208 : data_o = 1'b1;
            1209 : data_o = 1'b1;
            1210 : data_o = 1'b0;
            1211 : data_o = 1'b0;
            1212 : data_o = 1'b0;
            1213 : data_o = 1'b0;
            1214 : data_o = 1'b0;
            1215 : data_o = 1'b0;
            1216 : data_o = 1'b0;
            1217 : data_o = 1'b0;
            1218 : data_o = 1'b0;
            1219 : data_o = 1'b0;
            1220 : data_o = 1'b0;
            1221 : data_o = 1'b0;
            1222 : data_o = 1'b0;
            1223 : data_o = 1'b0;
            1224 : data_o = 1'b0;
            1225 : data_o = 1'b0;
            1226 : data_o = 1'b0;
            1227 : data_o = 1'b1;
            1228 : data_o = 1'b0;
            1229 : data_o = 1'b0;
            1230 : data_o = 1'b0;
            1231 : data_o = 1'b0;
            1232 : data_o = 1'b0;
            1233 : data_o = 1'b0;
            1234 : data_o = 1'b0;
            1235 : data_o = 1'b0;
            1236 : data_o = 1'b0;
            1237 : data_o = 1'b0;
            1238 : data_o = 1'b0;
            1239 : data_o = 1'b0;
            1240 : data_o = 1'b0;
            1241 : data_o = 1'b0;
            1242 : data_o = 1'b0;
            1243 : data_o = 1'b0;
            1244 : data_o = 1'b0;
            1245 : data_o = 1'b0;
            1246 : data_o = 1'b0;
            1247 : data_o = 1'b0;
            1248 : data_o = 1'b0;
            1249 : data_o = 1'b0;
            1250 : data_o = 1'b0;
            1251 : data_o = 1'b0;
            1252 : data_o = 1'b0;
            1253 : data_o = 1'b1;
            1254 : data_o = 1'b1;
            1255 : data_o = 1'b1;
            1256 : data_o = 1'b1;
            1257 : data_o = 1'b1;
            1258 : data_o = 1'b1;
            1259 : data_o = 1'b1;
            1260 : data_o = 1'b1;
            1261 : data_o = 1'b1;
            1262 : data_o = 1'b1;
            1263 : data_o = 1'b1;
            1264 : data_o = 1'b1;
            1265 : data_o = 1'b1;
            1266 : data_o = 1'b1;
            1267 : data_o = 1'b1;
            1268 : data_o = 1'b0;
            1269 : data_o = 1'b0;
            1270 : data_o = 1'b0;
            1271 : data_o = 1'b0;
            1272 : data_o = 1'b0;
            1273 : data_o = 1'b0;
            1274 : data_o = 1'b0;
            1275 : data_o = 1'b0;
            1276 : data_o = 1'b0;
            1277 : data_o = 1'b0;
            1278 : data_o = 1'b0;
            1279 : data_o = 1'b0;
            1280 : data_o = 1'b0;
            1281 : data_o = 1'b0;
            1282 : data_o = 1'b1;
            1283 : data_o = 1'b1;
            1284 : data_o = 1'b1;
            1285 : data_o = 1'b1;
            1286 : data_o = 1'b1;
            1287 : data_o = 1'b1;
            1288 : data_o = 1'b1;
            1289 : data_o = 1'b1;
            1290 : data_o = 1'b1;
            1291 : data_o = 1'b1;
            1292 : data_o = 1'b1;
            1293 : data_o = 1'b1;
            1294 : data_o = 1'b1;
            1295 : data_o = 1'b1;
            1296 : data_o = 1'b1;
            1297 : data_o = 1'b0;
            1298 : data_o = 1'b0;
            1299 : data_o = 1'b0;
            1300 : data_o = 1'b0;
            1301 : data_o = 1'b0;
            1302 : data_o = 1'b0;
            1303 : data_o = 1'b0;
            1304 : data_o = 1'b0;
            1305 : data_o = 1'b0;
            1306 : data_o = 1'b0;
            1307 : data_o = 1'b0;
            1308 : data_o = 1'b0;
            1309 : data_o = 1'b0;
            1310 : data_o = 1'b0;
            1311 : data_o = 1'b0;
            1312 : data_o = 1'b1;
            1313 : data_o = 1'b1;
            1314 : data_o = 1'b1;
            1315 : data_o = 1'b1;
            1316 : data_o = 1'b1;
            1317 : data_o = 1'b1;
            1318 : data_o = 1'b1;
            1319 : data_o = 1'b1;
            1320 : data_o = 1'b1;
            1321 : data_o = 1'b1;
            1322 : data_o = 1'b1;
            1323 : data_o = 1'b1;
            1324 : data_o = 1'b1;
            1325 : data_o = 1'b1;
            1326 : data_o = 1'b0;
            1327 : data_o = 1'b0;
            1328 : data_o = 1'b0;
            1329 : data_o = 1'b0;
            1330 : data_o = 1'b1;
            1331 : data_o = 1'b1;
            1332 : data_o = 1'b1;
            1333 : data_o = 1'b1;
            1334 : data_o = 1'b0;
            1335 : data_o = 1'b0;
            1336 : data_o = 1'b0;
            1337 : data_o = 1'b0;
            1338 : data_o = 1'b0;
            1339 : data_o = 1'b0;
            1340 : data_o = 1'b0;
            1341 : data_o = 1'b0;
            1342 : data_o = 1'b0;
            1343 : data_o = 1'b0;
            1344 : data_o = 1'b0;
            1345 : data_o = 1'b0;
            1346 : data_o = 1'b0;
            1347 : data_o = 1'b0;
            1348 : data_o = 1'b0;
            1349 : data_o = 1'b0;
            1350 : data_o = 1'b1;
            1351 : data_o = 1'b1;
            1352 : data_o = 1'b0;
            1353 : data_o = 1'b0;
            1354 : data_o = 1'b0;
            1355 : data_o = 1'b0;
            1356 : data_o = 1'b0;
            1357 : data_o = 1'b0;
            1358 : data_o = 1'b0;
            1359 : data_o = 1'b0;
            1360 : data_o = 1'b0;
            1361 : data_o = 1'b0;
            1362 : data_o = 1'b0;
            1363 : data_o = 1'b0;
            1364 : data_o = 1'b0;
            1365 : data_o = 1'b0;
            1366 : data_o = 1'b0;
            1367 : data_o = 1'b0;
            1368 : data_o = 1'b0;
            1369 : data_o = 1'b0;
            1370 : data_o = 1'b0;
            1371 : data_o = 1'b0;
            1372 : data_o = 1'b0;
            1373 : data_o = 1'b0;
            1374 : data_o = 1'b0;
            1375 : data_o = 1'b0;
            1376 : data_o = 1'b1;
            1377 : data_o = 1'b1;
            1378 : data_o = 1'b1;
            1379 : data_o = 1'b1;
            1380 : data_o = 1'b1;
            1381 : data_o = 1'b1;
            1382 : data_o = 1'b1;
            1383 : data_o = 1'b1;
            1384 : data_o = 1'b1;
            1385 : data_o = 1'b1;
            1386 : data_o = 1'b1;
            1387 : data_o = 1'b1;
            1388 : data_o = 1'b1;
            1389 : data_o = 1'b1;
            1390 : data_o = 1'b1;
            1391 : data_o = 1'b1;
            1392 : data_o = 1'b0;
            1393 : data_o = 1'b0;
            1394 : data_o = 1'b0;
            1395 : data_o = 1'b0;
            1396 : data_o = 1'b0;
            1397 : data_o = 1'b0;
            1398 : data_o = 1'b0;
            1399 : data_o = 1'b0;
            1400 : data_o = 1'b0;
            1401 : data_o = 1'b0;
            1402 : data_o = 1'b0;
            1403 : data_o = 1'b0;
            1404 : data_o = 1'b0;
            1405 : data_o = 1'b0;
            1406 : data_o = 1'b1;
            1407 : data_o = 1'b1;
            1408 : data_o = 1'b1;
            1409 : data_o = 1'b1;
            1410 : data_o = 1'b1;
            1411 : data_o = 1'b1;
            1412 : data_o = 1'b1;
            1413 : data_o = 1'b1;
            1414 : data_o = 1'b1;
            1415 : data_o = 1'b1;
            1416 : data_o = 1'b1;
            1417 : data_o = 1'b1;
            1418 : data_o = 1'b1;
            1419 : data_o = 1'b1;
            1420 : data_o = 1'b1;
            1421 : data_o = 1'b1;
            1422 : data_o = 1'b1;
            1423 : data_o = 1'b0;
            1424 : data_o = 1'b0;
            1425 : data_o = 1'b0;
            1426 : data_o = 1'b0;
            1427 : data_o = 1'b0;
            1428 : data_o = 1'b0;
            1429 : data_o = 1'b0;
            1430 : data_o = 1'b0;
            1431 : data_o = 1'b0;
            1432 : data_o = 1'b0;
            1433 : data_o = 1'b0;
            1434 : data_o = 1'b0;
            1435 : data_o = 1'b0;
            1436 : data_o = 1'b0;
            1437 : data_o = 1'b1;
            1438 : data_o = 1'b1;
            1439 : data_o = 1'b1;
            1440 : data_o = 1'b1;
            1441 : data_o = 1'b1;
            1442 : data_o = 1'b1;
            1443 : data_o = 1'b1;
            1444 : data_o = 1'b1;
            1445 : data_o = 1'b1;
            1446 : data_o = 1'b1;
            1447 : data_o = 1'b1;
            1448 : data_o = 1'b1;
            1449 : data_o = 1'b1;
            1450 : data_o = 1'b1;
            1451 : data_o = 1'b1;
            1452 : data_o = 1'b1;
            1453 : data_o = 1'b1;
            1454 : data_o = 1'b1;
            1455 : data_o = 1'b1;
            1456 : data_o = 1'b1;
            1457 : data_o = 1'b1;
            1458 : data_o = 1'b0;
            1459 : data_o = 1'b0;
            1460 : data_o = 1'b0;
            1461 : data_o = 1'b0;
            1462 : data_o = 1'b0;
            1463 : data_o = 1'b0;
            1464 : data_o = 1'b0;
            1465 : data_o = 1'b0;
            1466 : data_o = 1'b0;
            1467 : data_o = 1'b0;
            1468 : data_o = 1'b0;
            1469 : data_o = 1'b0;
            1470 : data_o = 1'b0;
            1471 : data_o = 1'b0;
            1472 : data_o = 1'b0;
            1473 : data_o = 1'b0;
            1474 : data_o = 1'b0;
            1475 : data_o = 1'b0;
            1476 : data_o = 1'b0;
            1477 : data_o = 1'b0;
            1478 : data_o = 1'b0;
            1479 : data_o = 1'b0;
            1480 : data_o = 1'b0;
            1481 : data_o = 1'b0;
            1482 : data_o = 1'b0;
            1483 : data_o = 1'b0;
            1484 : data_o = 1'b0;
            1485 : data_o = 1'b0;
            1486 : data_o = 1'b0;
            1487 : data_o = 1'b0;
            1488 : data_o = 1'b0;
            1489 : data_o = 1'b0;
            1490 : data_o = 1'b0;
            1491 : data_o = 1'b0;
            1492 : data_o = 1'b0;
            1493 : data_o = 1'b0;
            1494 : data_o = 1'b0;
            1495 : data_o = 1'b0;
            1496 : data_o = 1'b0;
            1497 : data_o = 1'b0;
            1498 : data_o = 1'b0;
            1499 : data_o = 1'b1;
            1500 : data_o = 1'b1;
            1501 : data_o = 1'b1;
            1502 : data_o = 1'b1;
            1503 : data_o = 1'b1;
            1504 : data_o = 1'b1;
            1505 : data_o = 1'b1;
            1506 : data_o = 1'b1;
            1507 : data_o = 1'b1;
            1508 : data_o = 1'b1;
            1509 : data_o = 1'b1;
            1510 : data_o = 1'b1;
            1511 : data_o = 1'b1;
            1512 : data_o = 1'b1;
            1513 : data_o = 1'b1;
            1514 : data_o = 1'b1;
            1515 : data_o = 1'b1;
            1516 : data_o = 1'b1;
            1517 : data_o = 1'b0;
            1518 : data_o = 1'b0;
            1519 : data_o = 1'b0;
            1520 : data_o = 1'b0;
            1521 : data_o = 1'b0;
            1522 : data_o = 1'b1;
            1523 : data_o = 1'b1;
            1524 : data_o = 1'b1;
            1525 : data_o = 1'b1;
            1526 : data_o = 1'b1;
            1527 : data_o = 1'b0;
            1528 : data_o = 1'b0;
            1529 : data_o = 1'b0;
            1530 : data_o = 1'b1;
            1531 : data_o = 1'b1;
            1532 : data_o = 1'b1;
            1533 : data_o = 1'b1;
            1534 : data_o = 1'b1;
            1535 : data_o = 1'b1;
            1536 : data_o = 1'b1;
            1537 : data_o = 1'b1;
            1538 : data_o = 1'b1;
            1539 : data_o = 1'b1;
            1540 : data_o = 1'b1;
            1541 : data_o = 1'b1;
            1542 : data_o = 1'b1;
            1543 : data_o = 1'b1;
            1544 : data_o = 1'b1;
            1545 : data_o = 1'b1;
            1546 : data_o = 1'b1;
            1547 : data_o = 1'b1;
            1548 : data_o = 1'b1;
            1549 : data_o = 1'b1;
            1550 : data_o = 1'b1;
            1551 : data_o = 1'b0;
            1552 : data_o = 1'b0;
            1553 : data_o = 1'b0;
            1554 : data_o = 1'b0;
            1555 : data_o = 1'b0;
            1556 : data_o = 1'b0;
            1557 : data_o = 1'b0;
            1558 : data_o = 1'b0;
            1559 : data_o = 1'b0;
            1560 : data_o = 1'b0;
            1561 : data_o = 1'b1;
            1562 : data_o = 1'b1;
            1563 : data_o = 1'b1;
            1564 : data_o = 1'b1;
            1565 : data_o = 1'b1;
            1566 : data_o = 1'b1;
            1567 : data_o = 1'b1;
            1568 : data_o = 1'b0;
            1569 : data_o = 1'b0;
            1570 : data_o = 1'b1;
            1571 : data_o = 1'b1;
            1572 : data_o = 1'b1;
            1573 : data_o = 1'b1;
            1574 : data_o = 1'b1;
            1575 : data_o = 1'b1;
            1576 : data_o = 1'b1;
            1577 : data_o = 1'b1;
            1578 : data_o = 1'b1;
            1579 : data_o = 1'b1;
            1580 : data_o = 1'b0;
            1581 : data_o = 1'b0;
            1582 : data_o = 1'b0;
            1583 : data_o = 1'b0;
            1584 : data_o = 1'b0;
            1585 : data_o = 1'b0;
            1586 : data_o = 1'b0;
            1587 : data_o = 1'b0;
            1588 : data_o = 1'b0;
            1589 : data_o = 1'b0;
            1590 : data_o = 1'b0;
            1591 : data_o = 1'b0;
            1592 : data_o = 1'b0;
            1593 : data_o = 1'b0;
            1594 : data_o = 1'b0;
            1595 : data_o = 1'b0;
            1596 : data_o = 1'b0;
            1597 : data_o = 1'b0;
            1598 : data_o = 1'b0;
            1599 : data_o = 1'b1;
            1600 : data_o = 1'b1;
            1601 : data_o = 1'b0;
            1602 : data_o = 1'b0;
            1603 : data_o = 1'b0;
            1604 : data_o = 1'b0;
            1605 : data_o = 1'b0;
            1606 : data_o = 1'b0;
            1607 : data_o = 1'b0;
            1608 : data_o = 1'b0;
            1609 : data_o = 1'b0;
            1610 : data_o = 1'b0;
            1611 : data_o = 1'b0;
            1612 : data_o = 1'b0;
            1613 : data_o = 1'b0;
            1614 : data_o = 1'b0;
            1615 : data_o = 1'b0;
            1616 : data_o = 1'b0;
            1617 : data_o = 1'b0;
            1618 : data_o = 1'b0;
            1619 : data_o = 1'b0;
            1620 : data_o = 1'b0;
            1621 : data_o = 1'b0;
            1622 : data_o = 1'b1;
            1623 : data_o = 1'b1;
            1624 : data_o = 1'b1;
            1625 : data_o = 1'b1;
            1626 : data_o = 1'b1;
            1627 : data_o = 1'b1;
            1628 : data_o = 1'b1;
            1629 : data_o = 1'b1;
            1630 : data_o = 1'b1;
            1631 : data_o = 1'b1;
            1632 : data_o = 1'b1;
            1633 : data_o = 1'b0;
            1634 : data_o = 1'b0;
            1635 : data_o = 1'b1;
            1636 : data_o = 1'b1;
            1637 : data_o = 1'b0;
            1638 : data_o = 1'b0;
            1639 : data_o = 1'b0;
            1640 : data_o = 1'b0;
            1641 : data_o = 1'b0;
            1642 : data_o = 1'b1;
            1643 : data_o = 1'b1;
            1644 : data_o = 1'b1;
            1645 : data_o = 1'b1;
            1646 : data_o = 1'b1;
            1647 : data_o = 1'b1;
            1648 : data_o = 1'b1;
            1649 : data_o = 1'b1;
            1650 : data_o = 1'b1;
            1651 : data_o = 1'b1;
            1652 : data_o = 1'b1;
            1653 : data_o = 1'b1;
            1654 : data_o = 1'b1;
            1655 : data_o = 1'b1;
            1656 : data_o = 1'b1;
            1657 : data_o = 1'b1;
            1658 : data_o = 1'b1;
            1659 : data_o = 1'b1;
            1660 : data_o = 1'b1;
            1661 : data_o = 1'b1;
            1662 : data_o = 1'b1;
            1663 : data_o = 1'b1;
            1664 : data_o = 1'b1;
            1665 : data_o = 1'b1;
            1666 : data_o = 1'b1;
            1667 : data_o = 1'b1;
            1668 : data_o = 1'b1;
            1669 : data_o = 1'b1;
            1670 : data_o = 1'b1;
            1671 : data_o = 1'b1;
            1672 : data_o = 1'b1;
            1673 : data_o = 1'b1;
            1674 : data_o = 1'b1;
            1675 : data_o = 1'b1;
            1676 : data_o = 1'b1;
            1677 : data_o = 1'b1;
            1678 : data_o = 1'b1;
            1679 : data_o = 1'b1;
            1680 : data_o = 1'b1;
            1681 : data_o = 1'b1;
            1682 : data_o = 1'b1;
            1683 : data_o = 1'b1;
            1684 : data_o = 1'b1;
            1685 : data_o = 1'b1;
            1686 : data_o = 1'b1;
            1687 : data_o = 1'b1;
            1688 : data_o = 1'b1;
            1689 : data_o = 1'b1;
            1690 : data_o = 1'b1;
            1691 : data_o = 1'b1;
            1692 : data_o = 1'b0;
            1693 : data_o = 1'b0;
            1694 : data_o = 1'b0;
            1695 : data_o = 1'b0;
            1696 : data_o = 1'b0;
            1697 : data_o = 1'b0;
            1698 : data_o = 1'b0;
            1699 : data_o = 1'b0;
            1700 : data_o = 1'b0;
            1701 : data_o = 1'b0;
            1702 : data_o = 1'b0;
            1703 : data_o = 1'b0;
            1704 : data_o = 1'b0;
            1705 : data_o = 1'b0;
            1706 : data_o = 1'b0;
            1707 : data_o = 1'b1;
            1708 : data_o = 1'b1;
            1709 : data_o = 1'b0;
            1710 : data_o = 1'b0;
            1711 : data_o = 1'b0;
            1712 : data_o = 1'b0;
            1713 : data_o = 1'b0;
            1714 : data_o = 1'b0;
            1715 : data_o = 1'b1;
            1716 : data_o = 1'b0;
            1717 : data_o = 1'b0;
            1718 : data_o = 1'b0;
            1719 : data_o = 1'b1;
            1720 : data_o = 1'b1;
            1721 : data_o = 1'b1;
            1722 : data_o = 1'b1;
            1723 : data_o = 1'b0;
            1724 : data_o = 1'b1;
            1725 : data_o = 1'b1;
            1726 : data_o = 1'b1;
            1727 : data_o = 1'b1;
            1728 : data_o = 1'b1;
            1729 : data_o = 1'b1;
            1730 : data_o = 1'b1;
            1731 : data_o = 1'b1;
            1732 : data_o = 1'b0;
            1733 : data_o = 1'b0;
            1734 : data_o = 1'b0;
            1735 : data_o = 1'b0;
            1736 : data_o = 1'b0;
            1737 : data_o = 1'b0;
            1738 : data_o = 1'b0;
            1739 : data_o = 1'b0;
            1740 : data_o = 1'b1;
            1741 : data_o = 1'b1;
            1742 : data_o = 1'b1;
            1743 : data_o = 1'b0;
            1744 : data_o = 1'b0;
            1745 : data_o = 1'b0;
            1746 : data_o = 1'b0;
            1747 : data_o = 1'b0;
            1748 : data_o = 1'b0;
            1749 : data_o = 1'b0;
            1750 : data_o = 1'b0;
            1751 : data_o = 1'b0;
            1752 : data_o = 1'b0;
            1753 : data_o = 1'b0;
            1754 : data_o = 1'b1;
            1755 : data_o = 1'b1;
            1756 : data_o = 1'b0;
            1757 : data_o = 1'b0;
            1758 : data_o = 1'b0;
            1759 : data_o = 1'b0;
            1760 : data_o = 1'b0;
            1761 : data_o = 1'b0;
            1762 : data_o = 1'b0;
            1763 : data_o = 1'b0;
            1764 : data_o = 1'b0;
            1765 : data_o = 1'b0;
            1766 : data_o = 1'b0;
            1767 : data_o = 1'b0;
            1768 : data_o = 1'b0;
            1769 : data_o = 1'b0;
            1770 : data_o = 1'b0;
            1771 : data_o = 1'b0;
            1772 : data_o = 1'b0;
            1773 : data_o = 1'b0;
            1774 : data_o = 1'b0;
            1775 : data_o = 1'b0;
            1776 : data_o = 1'b0;
            1777 : data_o = 1'b1;
            1778 : data_o = 1'b1;
            1779 : data_o = 1'b1;
            1780 : data_o = 1'b1;
            1781 : data_o = 1'b1;
            1782 : data_o = 1'b1;
            1783 : data_o = 1'b1;
            1784 : data_o = 1'b1;
            1785 : data_o = 1'b1;
            1786 : data_o = 1'b1;
            1787 : data_o = 1'b1;
            1788 : data_o = 1'b1;
            1789 : data_o = 1'b1;
            1790 : data_o = 1'b1;
            1791 : data_o = 1'b1;
            1792 : data_o = 1'b1;
            1793 : data_o = 1'b1;
            1794 : data_o = 1'b1;
            1795 : data_o = 1'b1;
            1796 : data_o = 1'b1;
            1797 : data_o = 1'b1;
            1798 : data_o = 1'b1;
            1799 : data_o = 1'b1;
            1800 : data_o = 1'b1;
            1801 : data_o = 1'b1;
            1802 : data_o = 1'b1;
            1803 : data_o = 1'b1;
            1804 : data_o = 1'b1;
            1805 : data_o = 1'b1;
            1806 : data_o = 1'b1;
            1807 : data_o = 1'b1;
            1808 : data_o = 1'b1;
            1809 : data_o = 1'b1;
            1810 : data_o = 1'b1;
            1811 : data_o = 1'b1;
            1812 : data_o = 1'b1;
            1813 : data_o = 1'b1;
            1814 : data_o = 1'b1;
            1815 : data_o = 1'b1;
            1816 : data_o = 1'b1;
            1817 : data_o = 1'b1;
            1818 : data_o = 1'b1;
            1819 : data_o = 1'b1;
            1820 : data_o = 1'b1;
            1821 : data_o = 1'b1;
            1822 : data_o = 1'b1;
            1823 : data_o = 1'b1;
            1824 : data_o = 1'b0;
            1825 : data_o = 1'b1;
            1826 : data_o = 1'b1;
            1827 : data_o = 1'b1;
            1828 : data_o = 1'b0;
            1829 : data_o = 1'b1;
            1830 : data_o = 1'b1;
            1831 : data_o = 1'b1;
            1832 : data_o = 1'b1;
            1833 : data_o = 1'b1;
            1834 : data_o = 1'b0;
            1835 : data_o = 1'b0;
            1836 : data_o = 1'b0;
            1837 : data_o = 1'b1;
            1838 : data_o = 1'b1;
            1839 : data_o = 1'b1;
            1840 : data_o = 1'b1;
            1841 : data_o = 1'b1;
            1842 : data_o = 1'b1;
            1843 : data_o = 1'b1;
            1844 : data_o = 1'b1;
            1845 : data_o = 1'b1;
            1846 : data_o = 1'b1;
            1847 : data_o = 1'b1;
            1848 : data_o = 1'b1;
            1849 : data_o = 1'b1;
            1850 : data_o = 1'b1;
            1851 : data_o = 1'b1;
            1852 : data_o = 1'b1;
            1853 : data_o = 1'b1;
            1854 : data_o = 1'b1;
            1855 : data_o = 1'b1;
            1856 : data_o = 1'b0;
            1857 : data_o = 1'b0;
            1858 : data_o = 1'b0;
            1859 : data_o = 1'b0;
            1860 : data_o = 1'b0;
            1861 : data_o = 1'b0;
            1862 : data_o = 1'b0;
            1863 : data_o = 1'b0;
            1864 : data_o = 1'b0;
            1865 : data_o = 1'b0;
            1866 : data_o = 1'b0;
            1867 : data_o = 1'b0;
            1868 : data_o = 1'b0;
            1869 : data_o = 1'b0;
            1870 : data_o = 1'b0;
            1871 : data_o = 1'b0;
            1872 : data_o = 1'b0;
            1873 : data_o = 1'b0;
            1874 : data_o = 1'b0;
            1875 : data_o = 1'b0;
            1876 : data_o = 1'b0;
            1877 : data_o = 1'b0;
            1878 : data_o = 1'b0;
            1879 : data_o = 1'b0;
            1880 : data_o = 1'b0;
            1881 : data_o = 1'b0;
            1882 : data_o = 1'b0;
            1883 : data_o = 1'b0;
            1884 : data_o = 1'b0;
            1885 : data_o = 1'b0;
            1886 : data_o = 1'b1;
            1887 : data_o = 1'b1;
            1888 : data_o = 1'b1;
            1889 : data_o = 1'b1;
            1890 : data_o = 1'b1;
            1891 : data_o = 1'b1;
            1892 : data_o = 1'b1;
            1893 : data_o = 1'b1;
            1894 : data_o = 1'b1;
            1895 : data_o = 1'b1;
            1896 : data_o = 1'b1;
            1897 : data_o = 1'b1;
            1898 : data_o = 1'b1;
            1899 : data_o = 1'b1;
            1900 : data_o = 1'b1;
            1901 : data_o = 1'b1;
            1902 : data_o = 1'b1;
            1903 : data_o = 1'b1;
            1904 : data_o = 1'b0;
            1905 : data_o = 1'b0;
            1906 : data_o = 1'b0;
            1907 : data_o = 1'b0;
            1908 : data_o = 1'b0;
            1909 : data_o = 1'b1;
            1910 : data_o = 1'b1;
            1911 : data_o = 1'b1;
            1912 : data_o = 1'b1;
            1913 : data_o = 1'b1;
            1914 : data_o = 1'b1;
            1915 : data_o = 1'b1;
            1916 : data_o = 1'b1;
            1917 : data_o = 1'b1;
            1918 : data_o = 1'b1;
            1919 : data_o = 1'b1;
            1920 : data_o = 1'b1;
            1921 : data_o = 1'b1;
            1922 : data_o = 1'b1;
            1923 : data_o = 1'b1;
            1924 : data_o = 1'b1;
            1925 : data_o = 1'b1;
            1926 : data_o = 1'b1;
            1927 : data_o = 1'b0;
            1928 : data_o = 1'b0;
            1929 : data_o = 1'b0;
            1930 : data_o = 1'b0;
            1931 : data_o = 1'b0;
            1932 : data_o = 1'b0;
            1933 : data_o = 1'b0;
            1934 : data_o = 1'b0;
            1935 : data_o = 1'b0;
            1936 : data_o = 1'b0;
            1937 : data_o = 1'b0;
            1938 : data_o = 1'b0;
            1939 : data_o = 1'b0;
            1940 : data_o = 1'b1;
            1941 : data_o = 1'b1;
            1942 : data_o = 1'b1;
            1943 : data_o = 1'b1;
            1944 : data_o = 1'b1;
            1945 : data_o = 1'b1;
            1946 : data_o = 1'b1;
            1947 : data_o = 1'b1;
            1948 : data_o = 1'b1;
            1949 : data_o = 1'b1;
            1950 : data_o = 1'b1;
            1951 : data_o = 1'b1;
            1952 : data_o = 1'b1;
            1953 : data_o = 1'b1;
            1954 : data_o = 1'b1;
            1955 : data_o = 1'b1;
            1956 : data_o = 1'b1;
            1957 : data_o = 1'b1;
            1958 : data_o = 1'b1;
            1959 : data_o = 1'b1;
            1960 : data_o = 1'b1;
            1961 : data_o = 1'b1;
            1962 : data_o = 1'b1;
            1963 : data_o = 1'b0;
            1964 : data_o = 1'b0;
            1965 : data_o = 1'b0;
            1966 : data_o = 1'b0;
            1967 : data_o = 1'b0;
            1968 : data_o = 1'b0;
            1969 : data_o = 1'b0;
            1970 : data_o = 1'b0;
            1971 : data_o = 1'b0;
            1972 : data_o = 1'b0;
            1973 : data_o = 1'b0;
            1974 : data_o = 1'b0;
            1975 : data_o = 1'b0;
            1976 : data_o = 1'b0;
            1977 : data_o = 1'b0;
            1978 : data_o = 1'b0;
            1979 : data_o = 1'b0;
            1980 : data_o = 1'b0;
            1981 : data_o = 1'b0;
            1982 : data_o = 1'b0;
            1983 : data_o = 1'b0;
            1984 : data_o = 1'b0;
            1985 : data_o = 1'b0;
            1986 : data_o = 1'b0;
            1987 : data_o = 1'b0;
            1988 : data_o = 1'b0;
            1989 : data_o = 1'b0;
            1990 : data_o = 1'b0;
            1991 : data_o = 1'b0;
            1992 : data_o = 1'b0;
            1993 : data_o = 1'b0;
            1994 : data_o = 1'b0;
            1995 : data_o = 1'b0;
            1996 : data_o = 1'b0;
            1997 : data_o = 1'b0;
            1998 : data_o = 1'b0;
            1999 : data_o = 1'b1;
            2000 : data_o = 1'b1;
            2001 : data_o = 1'b1;
            2002 : data_o = 1'b1;
            2003 : data_o = 1'b1;
            2004 : data_o = 1'b1;
            2005 : data_o = 1'b1;
            2006 : data_o = 1'b1;
            2007 : data_o = 1'b1;
            2008 : data_o = 1'b1;
            2009 : data_o = 1'b1;
            2010 : data_o = 1'b1;
            2011 : data_o = 1'b1;
            2012 : data_o = 1'b1;
            2013 : data_o = 1'b1;
            2014 : data_o = 1'b1;
            2015 : data_o = 1'b1;
            2016 : data_o = 1'b0;
            2017 : data_o = 1'b0;
            2018 : data_o = 1'b0;
            2019 : data_o = 1'b0;
            2020 : data_o = 1'b0;
            2021 : data_o = 1'b0;
            2022 : data_o = 1'b0;
            2023 : data_o = 1'b1;
            2024 : data_o = 1'b1;
            2025 : data_o = 1'b1;
            2026 : data_o = 1'b1;
            2027 : data_o = 1'b1;
            2028 : data_o = 1'b1;
            2029 : data_o = 1'b1;
            2030 : data_o = 1'b1;
            2031 : data_o = 1'b1;
            2032 : data_o = 1'b1;
            2033 : data_o = 1'b1;
            2034 : data_o = 1'b1;
            2035 : data_o = 1'b1;
            2036 : data_o = 1'b1;
            2037 : data_o = 1'b1;
            2038 : data_o = 1'b1;
            2039 : data_o = 1'b1;
            2040 : data_o = 1'b1;
            2041 : data_o = 1'b1;
            2042 : data_o = 1'b0;
            2043 : data_o = 1'b0;
            2044 : data_o = 1'b0;
            2045 : data_o = 1'b0;
            2046 : data_o = 1'b0;
            2047 : data_o = 1'b0;
            2048 : data_o = 1'b0;
            2049 : data_o = 1'b0;
            2050 : data_o = 1'b0;
            2051 : data_o = 1'b0;
            2052 : data_o = 1'b0;
            2053 : data_o = 1'b1;
            2054 : data_o = 1'b1;
            2055 : data_o = 1'b1;
            2056 : data_o = 1'b1;
            2057 : data_o = 1'b1;
            2058 : data_o = 1'b1;
            2059 : data_o = 1'b1;
            2060 : data_o = 1'b1;
            2061 : data_o = 1'b1;
            2062 : data_o = 1'b1;
            2063 : data_o = 1'b1;
            2064 : data_o = 1'b1;
            2065 : data_o = 1'b1;
            2066 : data_o = 1'b1;
            2067 : data_o = 1'b1;
            2068 : data_o = 1'b1;
            2069 : data_o = 1'b1;
            2070 : data_o = 1'b1;
            2071 : data_o = 1'b1;
            2072 : data_o = 1'b1;
            2073 : data_o = 1'b1;
            2074 : data_o = 1'b1;
            2075 : data_o = 1'b1;
            2076 : data_o = 1'b1;
            2077 : data_o = 1'b0;
            2078 : data_o = 1'b0;
            2079 : data_o = 1'b0;
            2080 : data_o = 1'b0;
            2081 : data_o = 1'b0;
            2082 : data_o = 1'b0;
            2083 : data_o = 1'b0;
            2084 : data_o = 1'b0;
            2085 : data_o = 1'b0;
            2086 : data_o = 1'b0;
            2087 : data_o = 1'b0;
            2088 : data_o = 1'b0;
            2089 : data_o = 1'b0;
            2090 : data_o = 1'b0;
            2091 : data_o = 1'b0;
            2092 : data_o = 1'b0;
            2093 : data_o = 1'b0;
            2094 : data_o = 1'b0;
            2095 : data_o = 1'b0;
            2096 : data_o = 1'b0;
            2097 : data_o = 1'b0;
            2098 : data_o = 1'b0;
            2099 : data_o = 1'b0;
            2100 : data_o = 1'b0;
            2101 : data_o = 1'b0;
            2102 : data_o = 1'b0;
            2103 : data_o = 1'b0;
            2104 : data_o = 1'b0;
            2105 : data_o = 1'b0;
            2106 : data_o = 1'b0;
            2107 : data_o = 1'b0;
            2108 : data_o = 1'b0;
            2109 : data_o = 1'b0;
            2110 : data_o = 1'b0;
            2111 : data_o = 1'b0;
            2112 : data_o = 1'b1;
            2113 : data_o = 1'b1;
            2114 : data_o = 1'b1;
            2115 : data_o = 1'b1;
            2116 : data_o = 1'b1;
            2117 : data_o = 1'b1;
            2118 : data_o = 1'b1;
            2119 : data_o = 1'b1;
            2120 : data_o = 1'b1;
            2121 : data_o = 1'b1;
            2122 : data_o = 1'b1;
            2123 : data_o = 1'b1;
            2124 : data_o = 1'b1;
            2125 : data_o = 1'b1;
            2126 : data_o = 1'b1;
            2127 : data_o = 1'b1;
            2128 : data_o = 1'b0;
            2129 : data_o = 1'b0;
            2130 : data_o = 1'b0;
            2131 : data_o = 1'b0;
            2132 : data_o = 1'b0;
            2133 : data_o = 1'b0;
            2134 : data_o = 1'b0;
            2135 : data_o = 1'b0;
            2136 : data_o = 1'b1;
            2137 : data_o = 1'b1;
            2138 : data_o = 1'b1;
            2139 : data_o = 1'b1;
            2140 : data_o = 1'b1;
            2141 : data_o = 1'b1;
            2142 : data_o = 1'b1;
            2143 : data_o = 1'b1;
            2144 : data_o = 1'b1;
            2145 : data_o = 1'b1;
            2146 : data_o = 1'b1;
            2147 : data_o = 1'b1;
            2148 : data_o = 1'b1;
            2149 : data_o = 1'b1;
            2150 : data_o = 1'b1;
            2151 : data_o = 1'b1;
            2152 : data_o = 1'b1;
            2153 : data_o = 1'b0;
            2154 : data_o = 1'b0;
            2155 : data_o = 1'b0;
            2156 : data_o = 1'b0;
            2157 : data_o = 1'b0;
            2158 : data_o = 1'b0;
            2159 : data_o = 1'b0;
            2160 : data_o = 1'b0;
            2161 : data_o = 1'b0;
            2162 : data_o = 1'b0;
            2163 : data_o = 1'b1;
            2164 : data_o = 1'b1;
            2165 : data_o = 1'b1;
            2166 : data_o = 1'b1;
            2167 : data_o = 1'b1;
            2168 : data_o = 1'b1;
            2169 : data_o = 1'b1;
            2170 : data_o = 1'b1;
            2171 : data_o = 1'b1;
            2172 : data_o = 1'b1;
            2173 : data_o = 1'b1;
            2174 : data_o = 1'b1;
            2175 : data_o = 1'b1;
            2176 : data_o = 1'b1;
            2177 : data_o = 1'b1;
            2178 : data_o = 1'b1;
            2179 : data_o = 1'b1;
            2180 : data_o = 1'b1;
            2181 : data_o = 1'b1;
            2182 : data_o = 1'b1;
            2183 : data_o = 1'b1;
            2184 : data_o = 1'b1;
            2185 : data_o = 1'b1;
            2186 : data_o = 1'b1;
            2187 : data_o = 1'b1;
            2188 : data_o = 1'b1;
            2189 : data_o = 1'b0;
            2190 : data_o = 1'b0;
            2191 : data_o = 1'b0;
            2192 : data_o = 1'b0;
            2193 : data_o = 1'b0;
            2194 : data_o = 1'b0;
            2195 : data_o = 1'b0;
            2196 : data_o = 1'b0;
            2197 : data_o = 1'b0;
            2198 : data_o = 1'b0;
            2199 : data_o = 1'b0;
            2200 : data_o = 1'b0;
            2201 : data_o = 1'b0;
            2202 : data_o = 1'b0;
            2203 : data_o = 1'b0;
            2204 : data_o = 1'b0;
            2205 : data_o = 1'b0;
            2206 : data_o = 1'b0;
            2207 : data_o = 1'b0;
            2208 : data_o = 1'b0;
            2209 : data_o = 1'b0;
            2210 : data_o = 1'b0;
            2211 : data_o = 1'b0;
            2212 : data_o = 1'b0;
            2213 : data_o = 1'b0;
            2214 : data_o = 1'b0;
            2215 : data_o = 1'b0;
            2216 : data_o = 1'b0;
            2217 : data_o = 1'b0;
            2218 : data_o = 1'b0;
            2219 : data_o = 1'b0;
            2220 : data_o = 1'b0;
            2221 : data_o = 1'b0;
            2222 : data_o = 1'b0;
            2223 : data_o = 1'b1;
            2224 : data_o = 1'b1;
            2225 : data_o = 1'b1;
            2226 : data_o = 1'b1;
            2227 : data_o = 1'b1;
            2228 : data_o = 1'b1;
            2229 : data_o = 1'b1;
            2230 : data_o = 1'b1;
            2231 : data_o = 1'b1;
            2232 : data_o = 1'b1;
            2233 : data_o = 1'b1;
            2234 : data_o = 1'b1;
            2235 : data_o = 1'b1;
            2236 : data_o = 1'b1;
            2237 : data_o = 1'b1;
            2238 : data_o = 1'b1;
            2239 : data_o = 1'b1;
            2240 : data_o = 1'b1;
            2241 : data_o = 1'b1;
            2242 : data_o = 1'b1;
            2243 : data_o = 1'b0;
            2244 : data_o = 1'b0;
            2245 : data_o = 1'b0;
            2246 : data_o = 1'b0;
            2247 : data_o = 1'b0;
            2248 : data_o = 1'b1;
            2249 : data_o = 1'b1;
            2250 : data_o = 1'b1;
            2251 : data_o = 1'b1;
            2252 : data_o = 1'b1;
            2253 : data_o = 1'b1;
            2254 : data_o = 1'b1;
            2255 : data_o = 1'b1;
            2256 : data_o = 1'b1;
            2257 : data_o = 1'b1;
            2258 : data_o = 1'b1;
            2259 : data_o = 1'b1;
            2260 : data_o = 1'b1;
            2261 : data_o = 1'b1;
            2262 : data_o = 1'b1;
            2263 : data_o = 1'b1;
            2264 : data_o = 1'b1;
            2265 : data_o = 1'b1;
            2266 : data_o = 1'b1;
            2267 : data_o = 1'b1;
            2268 : data_o = 1'b1;
            2269 : data_o = 1'b0;
            2270 : data_o = 1'b0;
            2271 : data_o = 1'b0;
            2272 : data_o = 1'b0;
            2273 : data_o = 1'b0;
            2274 : data_o = 1'b0;
            2275 : data_o = 1'b0;
            2276 : data_o = 1'b0;
            2277 : data_o = 1'b1;
            2278 : data_o = 1'b1;
            2279 : data_o = 1'b1;
            2280 : data_o = 1'b1;
            2281 : data_o = 1'b1;
            2282 : data_o = 1'b1;
            2283 : data_o = 1'b1;
            2284 : data_o = 1'b1;
            2285 : data_o = 1'b1;
            2286 : data_o = 1'b1;
            2287 : data_o = 1'b1;
            2288 : data_o = 1'b1;
            2289 : data_o = 1'b1;
            2290 : data_o = 1'b1;
            2291 : data_o = 1'b1;
            2292 : data_o = 1'b1;
            2293 : data_o = 1'b1;
            2294 : data_o = 1'b1;
            2295 : data_o = 1'b1;
            2296 : data_o = 1'b1;
            2297 : data_o = 1'b1;
            2298 : data_o = 1'b0;
            2299 : data_o = 1'b0;
            2300 : data_o = 1'b0;
            2301 : data_o = 1'b0;
            2302 : data_o = 1'b0;
            2303 : data_o = 1'b0;
            2304 : data_o = 1'b0;
            2305 : data_o = 1'b0;
            2306 : data_o = 1'b0;
            2307 : data_o = 1'b0;
            2308 : data_o = 1'b0;
            2309 : data_o = 1'b0;
            2310 : data_o = 1'b0;
            2311 : data_o = 1'b0;
            2312 : data_o = 1'b0;
            2313 : data_o = 1'b0;
            2314 : data_o = 1'b0;
            2315 : data_o = 1'b0;
            2316 : data_o = 1'b0;
            2317 : data_o = 1'b0;
            2318 : data_o = 1'b0;
            2319 : data_o = 1'b0;
            2320 : data_o = 1'b0;
            2321 : data_o = 1'b0;
            2322 : data_o = 1'b0;
            2323 : data_o = 1'b0;
            2324 : data_o = 1'b0;
            2325 : data_o = 1'b0;
            2326 : data_o = 1'b0;
            2327 : data_o = 1'b0;
            2328 : data_o = 1'b0;
            2329 : data_o = 1'b0;
            2330 : data_o = 1'b0;
            2331 : data_o = 1'b0;
            2332 : data_o = 1'b1;
            2333 : data_o = 1'b1;
            2334 : data_o = 1'b1;
            2335 : data_o = 1'b1;
            2336 : data_o = 1'b1;
            2337 : data_o = 1'b1;
            2338 : data_o = 1'b1;
            2339 : data_o = 1'b1;
            2340 : data_o = 1'b1;
            2341 : data_o = 1'b1;
            2342 : data_o = 1'b1;
            2343 : data_o = 1'b1;
            2344 : data_o = 1'b1;
            2345 : data_o = 1'b1;
            2346 : data_o = 1'b1;
            2347 : data_o = 1'b1;
            2348 : data_o = 1'b1;
            2349 : data_o = 1'b1;
            2350 : data_o = 1'b1;
            2351 : data_o = 1'b0;
            2352 : data_o = 1'b0;
            2353 : data_o = 1'b0;
            2354 : data_o = 1'b0;
            2355 : data_o = 1'b0;
            2356 : data_o = 1'b1;
            2357 : data_o = 1'b1;
            2358 : data_o = 1'b1;
            2359 : data_o = 1'b1;
            2360 : data_o = 1'b1;
            2361 : data_o = 1'b1;
            2362 : data_o = 1'b1;
            2363 : data_o = 1'b1;
            2364 : data_o = 1'b1;
            2365 : data_o = 1'b1;
            2366 : data_o = 1'b1;
            2367 : data_o = 1'b1;
            2368 : data_o = 1'b1;
            2369 : data_o = 1'b1;
            2370 : data_o = 1'b1;
            2371 : data_o = 1'b1;
            2372 : data_o = 1'b1;
            2373 : data_o = 1'b1;
            2374 : data_o = 1'b0;
            2375 : data_o = 1'b0;
            2376 : data_o = 1'b0;
            2377 : data_o = 1'b0;
            2378 : data_o = 1'b0;
            2379 : data_o = 1'b0;
            2380 : data_o = 1'b0;
            2381 : data_o = 1'b0;
            2382 : data_o = 1'b0;
            2383 : data_o = 1'b0;
            2384 : data_o = 1'b1;
            2385 : data_o = 1'b1;
            2386 : data_o = 1'b1;
            2387 : data_o = 1'b1;
            2388 : data_o = 1'b1;
            2389 : data_o = 1'b1;
            2390 : data_o = 1'b1;
            2391 : data_o = 1'b1;
            2392 : data_o = 1'b1;
            2393 : data_o = 1'b1;
            2394 : data_o = 1'b1;
            2395 : data_o = 1'b1;
            2396 : data_o = 1'b0;
            2397 : data_o = 1'b1;
            2398 : data_o = 1'b1;
            2399 : data_o = 1'b1;
            2400 : data_o = 1'b1;
            2401 : data_o = 1'b1;
            2402 : data_o = 1'b1;
            2403 : data_o = 1'b1;
            2404 : data_o = 1'b1;
            2405 : data_o = 1'b0;
            2406 : data_o = 1'b0;
            2407 : data_o = 1'b0;
            2408 : data_o = 1'b0;
            2409 : data_o = 1'b0;
            2410 : data_o = 1'b0;
            2411 : data_o = 1'b0;
            2412 : data_o = 1'b0;
            2413 : data_o = 1'b0;
            2414 : data_o = 1'b0;
            2415 : data_o = 1'b0;
            2416 : data_o = 1'b0;
            2417 : data_o = 1'b0;
            2418 : data_o = 1'b0;
            2419 : data_o = 1'b0;
            2420 : data_o = 1'b0;
            2421 : data_o = 1'b0;
            2422 : data_o = 1'b0;
            2423 : data_o = 1'b0;
            2424 : data_o = 1'b0;
            2425 : data_o = 1'b0;
            2426 : data_o = 1'b0;
            2427 : data_o = 1'b0;
            2428 : data_o = 1'b0;
            2429 : data_o = 1'b0;
            2430 : data_o = 1'b0;
            2431 : data_o = 1'b0;
            2432 : data_o = 1'b0;
            2433 : data_o = 1'b0;
            2434 : data_o = 1'b0;
            2435 : data_o = 1'b0;
            2436 : data_o = 1'b0;
            2437 : data_o = 1'b1;
            2438 : data_o = 1'b1;
            2439 : data_o = 1'b1;
            2440 : data_o = 1'b1;
            2441 : data_o = 1'b1;
            2442 : data_o = 1'b1;
            2443 : data_o = 1'b1;
            2444 : data_o = 1'b1;
            2445 : data_o = 1'b1;
            2446 : data_o = 1'b1;
            2447 : data_o = 1'b0;
            2448 : data_o = 1'b0;
            2449 : data_o = 1'b0;
            2450 : data_o = 1'b0;
            2451 : data_o = 1'b0;
            2452 : data_o = 1'b1;
            2453 : data_o = 1'b1;
            2454 : data_o = 1'b1;
            2455 : data_o = 1'b1;
            2456 : data_o = 1'b1;
            2457 : data_o = 1'b0;
            2458 : data_o = 1'b0;
            2459 : data_o = 1'b0;
            2460 : data_o = 1'b0;
            2461 : data_o = 1'b1;
            2462 : data_o = 1'b1;
            2463 : data_o = 1'b1;
            2464 : data_o = 1'b1;
            2465 : data_o = 1'b1;
            2466 : data_o = 1'b1;
            2467 : data_o = 1'b1;
            2468 : data_o = 1'b1;
            2469 : data_o = 1'b1;
            2470 : data_o = 1'b1;
            2471 : data_o = 1'b1;
            2472 : data_o = 1'b1;
            2473 : data_o = 1'b0;
            2474 : data_o = 1'b0;
            2475 : data_o = 1'b0;
            2476 : data_o = 1'b0;
            2477 : data_o = 1'b0;
            2478 : data_o = 1'b0;
            2479 : data_o = 1'b0;
            2480 : data_o = 1'b1;
            2481 : data_o = 1'b1;
            2482 : data_o = 1'b1;
            2483 : data_o = 1'b1;
            2484 : data_o = 1'b1;
            2485 : data_o = 1'b1;
            2486 : data_o = 1'b0;
            2487 : data_o = 1'b0;
            2488 : data_o = 1'b1;
            2489 : data_o = 1'b1;
            2490 : data_o = 1'b1;
            2491 : data_o = 1'b1;
            2492 : data_o = 1'b1;
            2493 : data_o = 1'b1;
            2494 : data_o = 1'b1;
            2495 : data_o = 1'b1;
            2496 : data_o = 1'b1;
            2497 : data_o = 1'b1;
            2498 : data_o = 1'b1;
            2499 : data_o = 1'b1;
            2500 : data_o = 1'b1;
            2501 : data_o = 1'b1;
            2502 : data_o = 1'b1;
            2503 : data_o = 1'b1;
            2504 : data_o = 1'b1;
            2505 : data_o = 1'b1;
            2506 : data_o = 1'b1;
            2507 : data_o = 1'b1;
            2508 : data_o = 1'b1;
            2509 : data_o = 1'b0;
            2510 : data_o = 1'b0;
            2511 : data_o = 1'b0;
            2512 : data_o = 1'b0;
            2513 : data_o = 1'b0;
            2514 : data_o = 1'b0;
            2515 : data_o = 1'b0;
            2516 : data_o = 1'b0;
            2517 : data_o = 1'b0;
            2518 : data_o = 1'b0;
            2519 : data_o = 1'b0;
            2520 : data_o = 1'b0;
            2521 : data_o = 1'b0;
            2522 : data_o = 1'b0;
            2523 : data_o = 1'b0;
            2524 : data_o = 1'b0;
            2525 : data_o = 1'b0;
            2526 : data_o = 1'b0;
            2527 : data_o = 1'b0;
            2528 : data_o = 1'b0;
            2529 : data_o = 1'b0;
            2530 : data_o = 1'b0;
            2531 : data_o = 1'b0;
            2532 : data_o = 1'b0;
            2533 : data_o = 1'b0;
            2534 : data_o = 1'b0;
            2535 : data_o = 1'b0;
            2536 : data_o = 1'b0;
            2537 : data_o = 1'b0;
            2538 : data_o = 1'b0;
            2539 : data_o = 1'b0;
            2540 : data_o = 1'b1;
            2541 : data_o = 1'b1;
            2542 : data_o = 1'b1;
            2543 : data_o = 1'b1;
            2544 : data_o = 1'b1;
            2545 : data_o = 1'b1;
            2546 : data_o = 1'b1;
            2547 : data_o = 1'b1;
            2548 : data_o = 1'b1;
            2549 : data_o = 1'b1;
            2550 : data_o = 1'b0;
            2551 : data_o = 1'b0;
            2552 : data_o = 1'b0;
            2553 : data_o = 1'b0;
            2554 : data_o = 1'b0;
            2555 : data_o = 1'b0;
            2556 : data_o = 1'b0;
            2557 : data_o = 1'b0;
            2558 : data_o = 1'b1;
            2559 : data_o = 1'b1;
            2560 : data_o = 1'b1;
            2561 : data_o = 1'b1;
            2562 : data_o = 1'b1;
            2563 : data_o = 1'b1;
            2564 : data_o = 1'b0;
            2565 : data_o = 1'b1;
            2566 : data_o = 1'b1;
            2567 : data_o = 1'b1;
            2568 : data_o = 1'b1;
            2569 : data_o = 1'b1;
            2570 : data_o = 1'b1;
            2571 : data_o = 1'b1;
            2572 : data_o = 1'b1;
            2573 : data_o = 1'b1;
            2574 : data_o = 1'b1;
            2575 : data_o = 1'b1;
            2576 : data_o = 1'b1;
            2577 : data_o = 1'b0;
            2578 : data_o = 1'b0;
            2579 : data_o = 1'b0;
            2580 : data_o = 1'b0;
            2581 : data_o = 1'b0;
            2582 : data_o = 1'b0;
            2583 : data_o = 1'b0;
            2584 : data_o = 1'b0;
            2585 : data_o = 1'b0;
            2586 : data_o = 1'b1;
            2587 : data_o = 1'b1;
            2588 : data_o = 1'b1;
            2589 : data_o = 1'b1;
            2590 : data_o = 1'b1;
            2591 : data_o = 1'b0;
            2592 : data_o = 1'b0;
            2593 : data_o = 1'b0;
            2594 : data_o = 1'b0;
            2595 : data_o = 1'b1;
            2596 : data_o = 1'b1;
            2597 : data_o = 1'b1;
            2598 : data_o = 1'b1;
            2599 : data_o = 1'b1;
            2600 : data_o = 1'b1;
            2601 : data_o = 1'b1;
            2602 : data_o = 1'b1;
            2603 : data_o = 1'b1;
            2604 : data_o = 1'b1;
            2605 : data_o = 1'b1;
            2606 : data_o = 1'b0;
            2607 : data_o = 1'b0;
            2608 : data_o = 1'b0;
            2609 : data_o = 1'b1;
            2610 : data_o = 1'b1;
            2611 : data_o = 1'b1;
            2612 : data_o = 1'b1;
            2613 : data_o = 1'b1;
            2614 : data_o = 1'b1;
            2615 : data_o = 1'b1;
            2616 : data_o = 1'b1;
            2617 : data_o = 1'b0;
            2618 : data_o = 1'b0;
            2619 : data_o = 1'b0;
            2620 : data_o = 1'b0;
            2621 : data_o = 1'b0;
            2622 : data_o = 1'b0;
            2623 : data_o = 1'b0;
            2624 : data_o = 1'b0;
            2625 : data_o = 1'b0;
            2626 : data_o = 1'b0;
            2627 : data_o = 1'b0;
            2628 : data_o = 1'b0;
            2629 : data_o = 1'b0;
            2630 : data_o = 1'b0;
            2631 : data_o = 1'b0;
            2632 : data_o = 1'b0;
            2633 : data_o = 1'b0;
            2634 : data_o = 1'b0;
            2635 : data_o = 1'b0;
            2636 : data_o = 1'b0;
            2637 : data_o = 1'b0;
            2638 : data_o = 1'b0;
            2639 : data_o = 1'b0;
            2640 : data_o = 1'b0;
            2641 : data_o = 1'b0;
            2642 : data_o = 1'b0;
            2643 : data_o = 1'b0;
            2644 : data_o = 1'b0;
            2645 : data_o = 1'b1;
            2646 : data_o = 1'b1;
            2647 : data_o = 1'b1;
            2648 : data_o = 1'b1;
            2649 : data_o = 1'b1;
            2650 : data_o = 1'b1;
            2651 : data_o = 1'b1;
            2652 : data_o = 1'b1;
            2653 : data_o = 1'b1;
            2654 : data_o = 1'b1;
            2655 : data_o = 1'b0;
            2656 : data_o = 1'b0;
            2657 : data_o = 1'b0;
            2658 : data_o = 1'b0;
            2659 : data_o = 1'b0;
            2660 : data_o = 1'b0;
            2661 : data_o = 1'b0;
            2662 : data_o = 1'b0;
            2663 : data_o = 1'b1;
            2664 : data_o = 1'b1;
            2665 : data_o = 1'b1;
            2666 : data_o = 1'b1;
            2667 : data_o = 1'b1;
            2668 : data_o = 1'b1;
            2669 : data_o = 1'b1;
            2670 : data_o = 1'b1;
            2671 : data_o = 1'b1;
            2672 : data_o = 1'b1;
            2673 : data_o = 1'b1;
            2674 : data_o = 1'b1;
            2675 : data_o = 1'b1;
            2676 : data_o = 1'b1;
            2677 : data_o = 1'b1;
            2678 : data_o = 1'b1;
            2679 : data_o = 1'b1;
            2680 : data_o = 1'b1;
            2681 : data_o = 1'b1;
            2682 : data_o = 1'b0;
            2683 : data_o = 1'b0;
            2684 : data_o = 1'b0;
            2685 : data_o = 1'b0;
            2686 : data_o = 1'b0;
            2687 : data_o = 1'b0;
            2688 : data_o = 1'b0;
            2689 : data_o = 1'b0;
            2690 : data_o = 1'b0;
            2691 : data_o = 1'b1;
            2692 : data_o = 1'b1;
            2693 : data_o = 1'b1;
            2694 : data_o = 1'b1;
            2695 : data_o = 1'b1;
            2696 : data_o = 1'b1;
            2697 : data_o = 1'b1;
            2698 : data_o = 1'b1;
            2699 : data_o = 1'b1;
            2700 : data_o = 1'b1;
            2701 : data_o = 1'b1;
            2702 : data_o = 1'b1;
            2703 : data_o = 1'b1;
            2704 : data_o = 1'b1;
            2705 : data_o = 1'b1;
            2706 : data_o = 1'b1;
            2707 : data_o = 1'b1;
            2708 : data_o = 1'b1;
            2709 : data_o = 1'b1;
            2710 : data_o = 1'b1;
            2711 : data_o = 1'b1;
            2712 : data_o = 1'b1;
            2713 : data_o = 1'b0;
            2714 : data_o = 1'b0;
            2715 : data_o = 1'b0;
            2716 : data_o = 1'b1;
            2717 : data_o = 1'b1;
            2718 : data_o = 1'b1;
            2719 : data_o = 1'b1;
            2720 : data_o = 1'b1;
            2721 : data_o = 1'b1;
            2722 : data_o = 1'b0;
            2723 : data_o = 1'b0;
            2724 : data_o = 1'b0;
            2725 : data_o = 1'b0;
            2726 : data_o = 1'b0;
            2727 : data_o = 1'b0;
            2728 : data_o = 1'b0;
            2729 : data_o = 1'b0;
            2730 : data_o = 1'b0;
            2731 : data_o = 1'b0;
            2732 : data_o = 1'b0;
            2733 : data_o = 1'b0;
            2734 : data_o = 1'b0;
            2735 : data_o = 1'b0;
            2736 : data_o = 1'b0;
            2737 : data_o = 1'b0;
            2738 : data_o = 1'b0;
            2739 : data_o = 1'b0;
            2740 : data_o = 1'b0;
            2741 : data_o = 1'b0;
            2742 : data_o = 1'b0;
            2743 : data_o = 1'b0;
            2744 : data_o = 1'b0;
            2745 : data_o = 1'b0;
            2746 : data_o = 1'b0;
            2747 : data_o = 1'b0;
            2748 : data_o = 1'b0;
            2749 : data_o = 1'b1;
            2750 : data_o = 1'b1;
            2751 : data_o = 1'b1;
            2752 : data_o = 1'b1;
            2753 : data_o = 1'b1;
            2754 : data_o = 1'b1;
            2755 : data_o = 1'b1;
            2756 : data_o = 1'b1;
            2757 : data_o = 1'b1;
            2758 : data_o = 1'b1;
            2759 : data_o = 1'b0;
            2760 : data_o = 1'b0;
            2761 : data_o = 1'b0;
            2762 : data_o = 1'b0;
            2763 : data_o = 1'b0;
            2764 : data_o = 1'b0;
            2765 : data_o = 1'b0;
            2766 : data_o = 1'b0;
            2767 : data_o = 1'b1;
            2768 : data_o = 1'b1;
            2769 : data_o = 1'b1;
            2770 : data_o = 1'b1;
            2771 : data_o = 1'b1;
            2772 : data_o = 1'b1;
            2773 : data_o = 1'b1;
            2774 : data_o = 1'b1;
            2775 : data_o = 1'b1;
            2776 : data_o = 1'b1;
            2777 : data_o = 1'b1;
            2778 : data_o = 1'b1;
            2779 : data_o = 1'b1;
            2780 : data_o = 1'b1;
            2781 : data_o = 1'b1;
            2782 : data_o = 1'b1;
            2783 : data_o = 1'b1;
            2784 : data_o = 1'b1;
            2785 : data_o = 1'b1;
            2786 : data_o = 1'b1;
            2787 : data_o = 1'b1;
            2788 : data_o = 1'b0;
            2789 : data_o = 1'b0;
            2790 : data_o = 1'b0;
            2791 : data_o = 1'b0;
            2792 : data_o = 1'b0;
            2793 : data_o = 1'b0;
            2794 : data_o = 1'b0;
            2795 : data_o = 1'b0;
            2796 : data_o = 1'b0;
            2797 : data_o = 1'b1;
            2798 : data_o = 1'b1;
            2799 : data_o = 1'b1;
            2800 : data_o = 1'b1;
            2801 : data_o = 1'b1;
            2802 : data_o = 1'b1;
            2803 : data_o = 1'b1;
            2804 : data_o = 1'b1;
            2805 : data_o = 1'b1;
            2806 : data_o = 1'b1;
            2807 : data_o = 1'b1;
            2808 : data_o = 1'b0;
            2809 : data_o = 1'b0;
            2810 : data_o = 1'b1;
            2811 : data_o = 1'b1;
            2812 : data_o = 1'b1;
            2813 : data_o = 1'b1;
            2814 : data_o = 1'b1;
            2815 : data_o = 1'b1;
            2816 : data_o = 1'b1;
            2817 : data_o = 1'b1;
            2818 : data_o = 1'b1;
            2819 : data_o = 1'b1;
            2820 : data_o = 1'b1;
            2821 : data_o = 1'b1;
            2822 : data_o = 1'b1;
            2823 : data_o = 1'b1;
            2824 : data_o = 1'b0;
            2825 : data_o = 1'b0;
            2826 : data_o = 1'b0;
            2827 : data_o = 1'b0;
            2828 : data_o = 1'b0;
            2829 : data_o = 1'b0;
            2830 : data_o = 1'b0;
            2831 : data_o = 1'b0;
            2832 : data_o = 1'b0;
            2833 : data_o = 1'b0;
            2834 : data_o = 1'b0;
            2835 : data_o = 1'b0;
            2836 : data_o = 1'b0;
            2837 : data_o = 1'b0;
            2838 : data_o = 1'b0;
            2839 : data_o = 1'b0;
            2840 : data_o = 1'b0;
            2841 : data_o = 1'b0;
            2842 : data_o = 1'b0;
            2843 : data_o = 1'b0;
            2844 : data_o = 1'b0;
            2845 : data_o = 1'b0;
            2846 : data_o = 1'b0;
            2847 : data_o = 1'b0;
            2848 : data_o = 1'b0;
            2849 : data_o = 1'b0;
            2850 : data_o = 1'b0;
            2851 : data_o = 1'b0;
            2852 : data_o = 1'b1;
            2853 : data_o = 1'b1;
            2854 : data_o = 1'b1;
            2855 : data_o = 1'b1;
            2856 : data_o = 1'b1;
            2857 : data_o = 1'b1;
            2858 : data_o = 1'b1;
            2859 : data_o = 1'b1;
            2860 : data_o = 1'b1;
            2861 : data_o = 1'b1;
            2862 : data_o = 1'b1;
            2863 : data_o = 1'b0;
            2864 : data_o = 1'b0;
            2865 : data_o = 1'b0;
            2866 : data_o = 1'b0;
            2867 : data_o = 1'b0;
            2868 : data_o = 1'b0;
            2869 : data_o = 1'b0;
            2870 : data_o = 1'b0;
            2871 : data_o = 1'b1;
            2872 : data_o = 1'b1;
            2873 : data_o = 1'b1;
            2874 : data_o = 1'b1;
            2875 : data_o = 1'b1;
            2876 : data_o = 1'b1;
            2877 : data_o = 1'b1;
            2878 : data_o = 1'b1;
            2879 : data_o = 1'b1;
            2880 : data_o = 1'b1;
            2881 : data_o = 1'b1;
            2882 : data_o = 1'b1;
            2883 : data_o = 1'b1;
            2884 : data_o = 1'b1;
            2885 : data_o = 1'b1;
            2886 : data_o = 1'b1;
            2887 : data_o = 1'b1;
            2888 : data_o = 1'b1;
            2889 : data_o = 1'b1;
            2890 : data_o = 1'b1;
            2891 : data_o = 1'b1;
            2892 : data_o = 1'b0;
            2893 : data_o = 1'b0;
            2894 : data_o = 1'b0;
            2895 : data_o = 1'b0;
            2896 : data_o = 1'b0;
            2897 : data_o = 1'b0;
            2898 : data_o = 1'b0;
            2899 : data_o = 1'b0;
            2900 : data_o = 1'b0;
            2901 : data_o = 1'b1;
            2902 : data_o = 1'b1;
            2903 : data_o = 1'b1;
            2904 : data_o = 1'b1;
            2905 : data_o = 1'b1;
            2906 : data_o = 1'b1;
            2907 : data_o = 1'b1;
            2908 : data_o = 1'b1;
            2909 : data_o = 1'b1;
            2910 : data_o = 1'b1;
            2911 : data_o = 1'b1;
            2912 : data_o = 1'b0;
            2913 : data_o = 1'b0;
            2914 : data_o = 1'b0;
            2915 : data_o = 1'b0;
            2916 : data_o = 1'b1;
            2917 : data_o = 1'b1;
            2918 : data_o = 1'b1;
            2919 : data_o = 1'b1;
            2920 : data_o = 1'b1;
            2921 : data_o = 1'b1;
            2922 : data_o = 1'b1;
            2923 : data_o = 1'b1;
            2924 : data_o = 1'b1;
            2925 : data_o = 1'b1;
            2926 : data_o = 1'b0;
            2927 : data_o = 1'b0;
            2928 : data_o = 1'b0;
            2929 : data_o = 1'b0;
            2930 : data_o = 1'b0;
            2931 : data_o = 1'b0;
            2932 : data_o = 1'b0;
            2933 : data_o = 1'b0;
            2934 : data_o = 1'b0;
            2935 : data_o = 1'b0;
            2936 : data_o = 1'b0;
            2937 : data_o = 1'b0;
            2938 : data_o = 1'b0;
            2939 : data_o = 1'b0;
            2940 : data_o = 1'b0;
            2941 : data_o = 1'b0;
            2942 : data_o = 1'b0;
            2943 : data_o = 1'b0;
            2944 : data_o = 1'b0;
            2945 : data_o = 1'b0;
            2946 : data_o = 1'b0;
            2947 : data_o = 1'b0;
            2948 : data_o = 1'b0;
            2949 : data_o = 1'b0;
            2950 : data_o = 1'b0;
            2951 : data_o = 1'b0;
            2952 : data_o = 1'b0;
            2953 : data_o = 1'b0;
            2954 : data_o = 1'b0;
            2955 : data_o = 1'b0;
            2956 : data_o = 1'b0;
            2957 : data_o = 1'b0;
            2958 : data_o = 1'b1;
            2959 : data_o = 1'b1;
            2960 : data_o = 1'b1;
            2961 : data_o = 1'b1;
            2962 : data_o = 1'b1;
            2963 : data_o = 1'b1;
            2964 : data_o = 1'b1;
            2965 : data_o = 1'b1;
            2966 : data_o = 1'b1;
            2967 : data_o = 1'b1;
            2968 : data_o = 1'b0;
            2969 : data_o = 1'b0;
            2970 : data_o = 1'b0;
            2971 : data_o = 1'b0;
            2972 : data_o = 1'b0;
            2973 : data_o = 1'b0;
            2974 : data_o = 1'b0;
            2975 : data_o = 1'b0;
            2976 : data_o = 1'b0;
            2977 : data_o = 1'b1;
            2978 : data_o = 1'b1;
            2979 : data_o = 1'b1;
            2980 : data_o = 1'b1;
            2981 : data_o = 1'b1;
            2982 : data_o = 1'b1;
            2983 : data_o = 1'b1;
            2984 : data_o = 1'b1;
            2985 : data_o = 1'b1;
            2986 : data_o = 1'b1;
            2987 : data_o = 1'b1;
            2988 : data_o = 1'b1;
            2989 : data_o = 1'b1;
            2990 : data_o = 1'b1;
            2991 : data_o = 1'b1;
            2992 : data_o = 1'b1;
            2993 : data_o = 1'b1;
            2994 : data_o = 1'b1;
            2995 : data_o = 1'b1;
            2996 : data_o = 1'b1;
            2997 : data_o = 1'b1;
            2998 : data_o = 1'b0;
            2999 : data_o = 1'b0;
            3000 : data_o = 1'b0;
            3001 : data_o = 1'b0;
            3002 : data_o = 1'b0;
            3003 : data_o = 1'b0;
            3004 : data_o = 1'b0;
            3005 : data_o = 1'b0;
            3006 : data_o = 1'b0;
            3007 : data_o = 1'b1;
            3008 : data_o = 1'b1;
            3009 : data_o = 1'b1;
            3010 : data_o = 1'b1;
            3011 : data_o = 1'b1;
            3012 : data_o = 1'b1;
            3013 : data_o = 1'b1;
            3014 : data_o = 1'b1;
            3015 : data_o = 1'b1;
            3016 : data_o = 1'b1;
            3017 : data_o = 1'b1;
            3018 : data_o = 1'b0;
            3019 : data_o = 1'b0;
            3020 : data_o = 1'b0;
            3021 : data_o = 1'b0;
            3022 : data_o = 1'b0;
            3023 : data_o = 1'b0;
            3024 : data_o = 1'b1;
            3025 : data_o = 1'b1;
            3026 : data_o = 1'b1;
            3027 : data_o = 1'b1;
            3028 : data_o = 1'b1;
            3029 : data_o = 1'b1;
            3030 : data_o = 1'b1;
            3031 : data_o = 1'b1;
            3032 : data_o = 1'b1;
            3033 : data_o = 1'b0;
            3034 : data_o = 1'b0;
            3035 : data_o = 1'b0;
            3036 : data_o = 1'b0;
            3037 : data_o = 1'b0;
            3038 : data_o = 1'b0;
            3039 : data_o = 1'b0;
            3040 : data_o = 1'b0;
            3041 : data_o = 1'b0;
            3042 : data_o = 1'b0;
            3043 : data_o = 1'b0;
            3044 : data_o = 1'b0;
            3045 : data_o = 1'b0;
            3046 : data_o = 1'b0;
            3047 : data_o = 1'b0;
            3048 : data_o = 1'b0;
            3049 : data_o = 1'b0;
            3050 : data_o = 1'b0;
            3051 : data_o = 1'b0;
            3052 : data_o = 1'b0;
            3053 : data_o = 1'b0;
            3054 : data_o = 1'b0;
            3055 : data_o = 1'b0;
            3056 : data_o = 1'b0;
            3057 : data_o = 1'b0;
            3058 : data_o = 1'b0;
            3059 : data_o = 1'b0;
            3060 : data_o = 1'b0;
            3061 : data_o = 1'b0;
            3062 : data_o = 1'b1;
            3063 : data_o = 1'b1;
            3064 : data_o = 1'b1;
            3065 : data_o = 1'b1;
            3066 : data_o = 1'b1;
            3067 : data_o = 1'b1;
            3068 : data_o = 1'b1;
            3069 : data_o = 1'b1;
            3070 : data_o = 1'b1;
            3071 : data_o = 1'b1;
            3072 : data_o = 1'b1;
            3073 : data_o = 1'b0;
            3074 : data_o = 1'b0;
            3075 : data_o = 1'b0;
            3076 : data_o = 1'b0;
            3077 : data_o = 1'b0;
            3078 : data_o = 1'b0;
            3079 : data_o = 1'b0;
            3080 : data_o = 1'b0;
            3081 : data_o = 1'b0;
            3082 : data_o = 1'b1;
            3083 : data_o = 1'b1;
            3084 : data_o = 1'b1;
            3085 : data_o = 1'b1;
            3086 : data_o = 1'b1;
            3087 : data_o = 1'b1;
            3088 : data_o = 1'b1;
            3089 : data_o = 1'b1;
            3090 : data_o = 1'b1;
            3091 : data_o = 1'b1;
            3092 : data_o = 1'b1;
            3093 : data_o = 1'b1;
            3094 : data_o = 1'b1;
            3095 : data_o = 1'b1;
            3096 : data_o = 1'b1;
            3097 : data_o = 1'b1;
            3098 : data_o = 1'b1;
            3099 : data_o = 1'b1;
            3100 : data_o = 1'b1;
            3101 : data_o = 1'b1;
            3102 : data_o = 1'b1;
            3103 : data_o = 1'b1;
            3104 : data_o = 1'b1;
            3105 : data_o = 1'b0;
            3106 : data_o = 1'b0;
            3107 : data_o = 1'b0;
            3108 : data_o = 1'b0;
            3109 : data_o = 1'b0;
            3110 : data_o = 1'b0;
            3111 : data_o = 1'b0;
            3112 : data_o = 1'b0;
            3113 : data_o = 1'b0;
            3114 : data_o = 1'b0;
            3115 : data_o = 1'b1;
            3116 : data_o = 1'b1;
            3117 : data_o = 1'b1;
            3118 : data_o = 1'b1;
            3119 : data_o = 1'b1;
            3120 : data_o = 1'b1;
            3121 : data_o = 1'b1;
            3122 : data_o = 1'b1;
            3123 : data_o = 1'b1;
            3124 : data_o = 1'b1;
            3125 : data_o = 1'b0;
            3126 : data_o = 1'b0;
            3127 : data_o = 1'b0;
            3128 : data_o = 1'b0;
            3129 : data_o = 1'b0;
            3130 : data_o = 1'b0;
            3131 : data_o = 1'b0;
            3132 : data_o = 1'b0;
            3133 : data_o = 1'b1;
            3134 : data_o = 1'b1;
            3135 : data_o = 1'b1;
            3136 : data_o = 1'b1;
            3137 : data_o = 1'b1;
            3138 : data_o = 1'b1;
            3139 : data_o = 1'b1;
            3140 : data_o = 1'b0;
            3141 : data_o = 1'b0;
            3142 : data_o = 1'b0;
            3143 : data_o = 1'b0;
            3144 : data_o = 1'b0;
            3145 : data_o = 1'b0;
            3146 : data_o = 1'b0;
            3147 : data_o = 1'b0;
            3148 : data_o = 1'b0;
            3149 : data_o = 1'b0;
            3150 : data_o = 1'b0;
            3151 : data_o = 1'b0;
            3152 : data_o = 1'b0;
            3153 : data_o = 1'b0;
            3154 : data_o = 1'b0;
            3155 : data_o = 1'b0;
            3156 : data_o = 1'b0;
            3157 : data_o = 1'b0;
            3158 : data_o = 1'b0;
            3159 : data_o = 1'b0;
            3160 : data_o = 1'b0;
            3161 : data_o = 1'b0;
            3162 : data_o = 1'b0;
            3163 : data_o = 1'b0;
            3164 : data_o = 1'b0;
            3165 : data_o = 1'b0;
            3166 : data_o = 1'b0;
            3167 : data_o = 1'b0;
            3168 : data_o = 1'b1;
            3169 : data_o = 1'b1;
            3170 : data_o = 1'b1;
            3171 : data_o = 1'b1;
            3172 : data_o = 1'b1;
            3173 : data_o = 1'b1;
            3174 : data_o = 1'b1;
            3175 : data_o = 1'b1;
            3176 : data_o = 1'b1;
            3177 : data_o = 1'b1;
            3178 : data_o = 1'b1;
            3179 : data_o = 1'b0;
            3180 : data_o = 1'b0;
            3181 : data_o = 1'b0;
            3182 : data_o = 1'b0;
            3183 : data_o = 1'b0;
            3184 : data_o = 1'b0;
            3185 : data_o = 1'b0;
            3186 : data_o = 1'b0;
            3187 : data_o = 1'b0;
            3188 : data_o = 1'b1;
            3189 : data_o = 1'b1;
            3190 : data_o = 1'b1;
            3191 : data_o = 1'b1;
            3192 : data_o = 1'b1;
            3193 : data_o = 1'b1;
            3194 : data_o = 1'b1;
            3195 : data_o = 1'b1;
            3196 : data_o = 1'b1;
            3197 : data_o = 1'b1;
            3198 : data_o = 1'b1;
            3199 : data_o = 1'b1;
            3200 : data_o = 1'b1;
            3201 : data_o = 1'b0;
            3202 : data_o = 1'b0;
            3203 : data_o = 1'b1;
            3204 : data_o = 1'b1;
            3205 : data_o = 1'b1;
            3206 : data_o = 1'b1;
            3207 : data_o = 1'b1;
            3208 : data_o = 1'b1;
            3209 : data_o = 1'b1;
            3210 : data_o = 1'b1;
            3211 : data_o = 1'b1;
            3212 : data_o = 1'b1;
            3213 : data_o = 1'b0;
            3214 : data_o = 1'b0;
            3215 : data_o = 1'b0;
            3216 : data_o = 1'b0;
            3217 : data_o = 1'b0;
            3218 : data_o = 1'b0;
            3219 : data_o = 1'b0;
            3220 : data_o = 1'b0;
            3221 : data_o = 1'b1;
            3222 : data_o = 1'b1;
            3223 : data_o = 1'b1;
            3224 : data_o = 1'b1;
            3225 : data_o = 1'b1;
            3226 : data_o = 1'b1;
            3227 : data_o = 1'b1;
            3228 : data_o = 1'b1;
            3229 : data_o = 1'b1;
            3230 : data_o = 1'b1;
            3231 : data_o = 1'b0;
            3232 : data_o = 1'b0;
            3233 : data_o = 1'b0;
            3234 : data_o = 1'b0;
            3235 : data_o = 1'b0;
            3236 : data_o = 1'b0;
            3237 : data_o = 1'b0;
            3238 : data_o = 1'b0;
            3239 : data_o = 1'b0;
            3240 : data_o = 1'b1;
            3241 : data_o = 1'b1;
            3242 : data_o = 1'b1;
            3243 : data_o = 1'b1;
            3244 : data_o = 1'b1;
            3245 : data_o = 1'b0;
            3246 : data_o = 1'b0;
            3247 : data_o = 1'b0;
            3248 : data_o = 1'b0;
            3249 : data_o = 1'b0;
            3250 : data_o = 1'b0;
            3251 : data_o = 1'b0;
            3252 : data_o = 1'b0;
            3253 : data_o = 1'b0;
            3254 : data_o = 1'b0;
            3255 : data_o = 1'b0;
            3256 : data_o = 1'b0;
            3257 : data_o = 1'b0;
            3258 : data_o = 1'b0;
            3259 : data_o = 1'b0;
            3260 : data_o = 1'b0;
            3261 : data_o = 1'b0;
            3262 : data_o = 1'b0;
            3263 : data_o = 1'b0;
            3264 : data_o = 1'b0;
            3265 : data_o = 1'b0;
            3266 : data_o = 1'b0;
            3267 : data_o = 1'b0;
            3268 : data_o = 1'b0;
            3269 : data_o = 1'b0;
            3270 : data_o = 1'b0;
            3271 : data_o = 1'b0;
            3272 : data_o = 1'b1;
            3273 : data_o = 1'b1;
            3274 : data_o = 1'b1;
            3275 : data_o = 1'b1;
            3276 : data_o = 1'b1;
            3277 : data_o = 1'b1;
            3278 : data_o = 1'b1;
            3279 : data_o = 1'b1;
            3280 : data_o = 1'b1;
            3281 : data_o = 1'b1;
            3282 : data_o = 1'b1;
            3283 : data_o = 1'b0;
            3284 : data_o = 1'b0;
            3285 : data_o = 1'b0;
            3286 : data_o = 1'b0;
            3287 : data_o = 1'b0;
            3288 : data_o = 1'b0;
            3289 : data_o = 1'b0;
            3290 : data_o = 1'b0;
            3291 : data_o = 1'b0;
            3292 : data_o = 1'b0;
            3293 : data_o = 1'b1;
            3294 : data_o = 1'b1;
            3295 : data_o = 1'b1;
            3296 : data_o = 1'b1;
            3297 : data_o = 1'b1;
            3298 : data_o = 1'b1;
            3299 : data_o = 1'b1;
            3300 : data_o = 1'b1;
            3301 : data_o = 1'b1;
            3302 : data_o = 1'b1;
            3303 : data_o = 1'b1;
            3304 : data_o = 1'b1;
            3305 : data_o = 1'b0;
            3306 : data_o = 1'b0;
            3307 : data_o = 1'b0;
            3308 : data_o = 1'b0;
            3309 : data_o = 1'b0;
            3310 : data_o = 1'b0;
            3311 : data_o = 1'b0;
            3312 : data_o = 1'b1;
            3313 : data_o = 1'b1;
            3314 : data_o = 1'b1;
            3315 : data_o = 1'b1;
            3316 : data_o = 1'b1;
            3317 : data_o = 1'b1;
            3318 : data_o = 1'b1;
            3319 : data_o = 1'b1;
            3320 : data_o = 1'b1;
            3321 : data_o = 1'b1;
            3322 : data_o = 1'b0;
            3323 : data_o = 1'b0;
            3324 : data_o = 1'b0;
            3325 : data_o = 1'b0;
            3326 : data_o = 1'b0;
            3327 : data_o = 1'b1;
            3328 : data_o = 1'b1;
            3329 : data_o = 1'b1;
            3330 : data_o = 1'b1;
            3331 : data_o = 1'b1;
            3332 : data_o = 1'b1;
            3333 : data_o = 1'b1;
            3334 : data_o = 1'b1;
            3335 : data_o = 1'b1;
            3336 : data_o = 1'b1;
            3337 : data_o = 1'b1;
            3338 : data_o = 1'b1;
            3339 : data_o = 1'b1;
            3340 : data_o = 1'b1;
            3341 : data_o = 1'b1;
            3342 : data_o = 1'b0;
            3343 : data_o = 1'b0;
            3344 : data_o = 1'b0;
            3345 : data_o = 1'b0;
            3346 : data_o = 1'b0;
            3347 : data_o = 1'b0;
            3348 : data_o = 1'b0;
            3349 : data_o = 1'b0;
            3350 : data_o = 1'b0;
            3351 : data_o = 1'b0;
            3352 : data_o = 1'b0;
            3353 : data_o = 1'b0;
            3354 : data_o = 1'b0;
            3355 : data_o = 1'b0;
            3356 : data_o = 1'b0;
            3357 : data_o = 1'b0;
            3358 : data_o = 1'b0;
            3359 : data_o = 1'b0;
            3360 : data_o = 1'b0;
            3361 : data_o = 1'b0;
            3362 : data_o = 1'b0;
            3363 : data_o = 1'b0;
            3364 : data_o = 1'b0;
            3365 : data_o = 1'b0;
            3366 : data_o = 1'b0;
            3367 : data_o = 1'b0;
            3368 : data_o = 1'b0;
            3369 : data_o = 1'b0;
            3370 : data_o = 1'b0;
            3371 : data_o = 1'b0;
            3372 : data_o = 1'b0;
            3373 : data_o = 1'b0;
            3374 : data_o = 1'b0;
            3375 : data_o = 1'b0;
            3376 : data_o = 1'b0;
            3377 : data_o = 1'b1;
            3378 : data_o = 1'b1;
            3379 : data_o = 1'b1;
            3380 : data_o = 1'b1;
            3381 : data_o = 1'b1;
            3382 : data_o = 1'b1;
            3383 : data_o = 1'b1;
            3384 : data_o = 1'b1;
            3385 : data_o = 1'b1;
            3386 : data_o = 1'b1;
            3387 : data_o = 1'b1;
            3388 : data_o = 1'b0;
            3389 : data_o = 1'b0;
            3390 : data_o = 1'b0;
            3391 : data_o = 1'b0;
            3392 : data_o = 1'b0;
            3393 : data_o = 1'b0;
            3394 : data_o = 1'b0;
            3395 : data_o = 1'b0;
            3396 : data_o = 1'b0;
            3397 : data_o = 1'b0;
            3398 : data_o = 1'b1;
            3399 : data_o = 1'b1;
            3400 : data_o = 1'b1;
            3401 : data_o = 1'b1;
            3402 : data_o = 1'b1;
            3403 : data_o = 1'b1;
            3404 : data_o = 1'b1;
            3405 : data_o = 1'b1;
            3406 : data_o = 1'b1;
            3407 : data_o = 1'b1;
            3408 : data_o = 1'b1;
            3409 : data_o = 1'b1;
            3410 : data_o = 1'b1;
            3411 : data_o = 1'b0;
            3412 : data_o = 1'b0;
            3413 : data_o = 1'b0;
            3414 : data_o = 1'b0;
            3415 : data_o = 1'b0;
            3416 : data_o = 1'b0;
            3417 : data_o = 1'b0;
            3418 : data_o = 1'b0;
            3419 : data_o = 1'b1;
            3420 : data_o = 1'b1;
            3421 : data_o = 1'b1;
            3422 : data_o = 1'b1;
            3423 : data_o = 1'b1;
            3424 : data_o = 1'b1;
            3425 : data_o = 1'b1;
            3426 : data_o = 1'b1;
            3427 : data_o = 1'b1;
            3428 : data_o = 1'b1;
            3429 : data_o = 1'b1;
            3430 : data_o = 1'b0;
            3431 : data_o = 1'b0;
            3432 : data_o = 1'b0;
            3433 : data_o = 1'b0;
            3434 : data_o = 1'b0;
            3435 : data_o = 1'b0;
            3436 : data_o = 1'b0;
            3437 : data_o = 1'b1;
            3438 : data_o = 1'b1;
            3439 : data_o = 1'b1;
            3440 : data_o = 1'b1;
            3441 : data_o = 1'b1;
            3442 : data_o = 1'b1;
            3443 : data_o = 1'b1;
            3444 : data_o = 1'b1;
            3445 : data_o = 1'b1;
            3446 : data_o = 1'b1;
            3447 : data_o = 1'b1;
            3448 : data_o = 1'b1;
            3449 : data_o = 1'b1;
            3450 : data_o = 1'b0;
            3451 : data_o = 1'b0;
            3452 : data_o = 1'b0;
            3453 : data_o = 1'b0;
            3454 : data_o = 1'b0;
            3455 : data_o = 1'b0;
            3456 : data_o = 1'b0;
            3457 : data_o = 1'b0;
            3458 : data_o = 1'b0;
            3459 : data_o = 1'b0;
            3460 : data_o = 1'b0;
            3461 : data_o = 1'b0;
            3462 : data_o = 1'b0;
            3463 : data_o = 1'b0;
            3464 : data_o = 1'b0;
            3465 : data_o = 1'b0;
            3466 : data_o = 1'b0;
            3467 : data_o = 1'b0;
            3468 : data_o = 1'b0;
            3469 : data_o = 1'b0;
            3470 : data_o = 1'b0;
            3471 : data_o = 1'b0;
            3472 : data_o = 1'b0;
            3473 : data_o = 1'b0;
            3474 : data_o = 1'b0;
            3475 : data_o = 1'b0;
            3476 : data_o = 1'b0;
            3477 : data_o = 1'b0;
            3478 : data_o = 1'b0;
            3479 : data_o = 1'b0;
            3480 : data_o = 1'b0;
            3481 : data_o = 1'b0;
            3482 : data_o = 1'b1;
            3483 : data_o = 1'b1;
            3484 : data_o = 1'b1;
            3485 : data_o = 1'b1;
            3486 : data_o = 1'b1;
            3487 : data_o = 1'b1;
            3488 : data_o = 1'b1;
            3489 : data_o = 1'b1;
            3490 : data_o = 1'b1;
            3491 : data_o = 1'b1;
            3492 : data_o = 1'b1;
            3493 : data_o = 1'b1;
            3494 : data_o = 1'b0;
            3495 : data_o = 1'b0;
            3496 : data_o = 1'b0;
            3497 : data_o = 1'b0;
            3498 : data_o = 1'b0;
            3499 : data_o = 1'b0;
            3500 : data_o = 1'b0;
            3501 : data_o = 1'b0;
            3502 : data_o = 1'b0;
            3503 : data_o = 1'b0;
            3504 : data_o = 1'b1;
            3505 : data_o = 1'b1;
            3506 : data_o = 1'b1;
            3507 : data_o = 1'b1;
            3508 : data_o = 1'b1;
            3509 : data_o = 1'b1;
            3510 : data_o = 1'b1;
            3511 : data_o = 1'b1;
            3512 : data_o = 1'b1;
            3513 : data_o = 1'b1;
            3514 : data_o = 1'b1;
            3515 : data_o = 1'b1;
            3516 : data_o = 1'b1;
            3517 : data_o = 1'b1;
            3518 : data_o = 1'b0;
            3519 : data_o = 1'b0;
            3520 : data_o = 1'b0;
            3521 : data_o = 1'b0;
            3522 : data_o = 1'b0;
            3523 : data_o = 1'b0;
            3524 : data_o = 1'b0;
            3525 : data_o = 1'b0;
            3526 : data_o = 1'b0;
            3527 : data_o = 1'b1;
            3528 : data_o = 1'b1;
            3529 : data_o = 1'b1;
            3530 : data_o = 1'b1;
            3531 : data_o = 1'b1;
            3532 : data_o = 1'b1;
            3533 : data_o = 1'b1;
            3534 : data_o = 1'b1;
            3535 : data_o = 1'b1;
            3536 : data_o = 1'b1;
            3537 : data_o = 1'b1;
            3538 : data_o = 1'b1;
            3539 : data_o = 1'b1;
            3540 : data_o = 1'b1;
            3541 : data_o = 1'b0;
            3542 : data_o = 1'b0;
            3543 : data_o = 1'b0;
            3544 : data_o = 1'b0;
            3545 : data_o = 1'b0;
            3546 : data_o = 1'b1;
            3547 : data_o = 1'b1;
            3548 : data_o = 1'b1;
            3549 : data_o = 1'b1;
            3550 : data_o = 1'b1;
            3551 : data_o = 1'b1;
            3552 : data_o = 1'b1;
            3553 : data_o = 1'b1;
            3554 : data_o = 1'b1;
            3555 : data_o = 1'b1;
            3556 : data_o = 1'b1;
            3557 : data_o = 1'b1;
            3558 : data_o = 1'b0;
            3559 : data_o = 1'b0;
            3560 : data_o = 1'b0;
            3561 : data_o = 1'b0;
            3562 : data_o = 1'b0;
            3563 : data_o = 1'b0;
            3564 : data_o = 1'b0;
            3565 : data_o = 1'b0;
            3566 : data_o = 1'b0;
            3567 : data_o = 1'b0;
            3568 : data_o = 1'b0;
            3569 : data_o = 1'b0;
            3570 : data_o = 1'b0;
            3571 : data_o = 1'b0;
            3572 : data_o = 1'b0;
            3573 : data_o = 1'b0;
            3574 : data_o = 1'b0;
            3575 : data_o = 1'b0;
            3576 : data_o = 1'b0;
            3577 : data_o = 1'b0;
            3578 : data_o = 1'b0;
            3579 : data_o = 1'b0;
            3580 : data_o = 1'b0;
            3581 : data_o = 1'b0;
            3582 : data_o = 1'b0;
            3583 : data_o = 1'b0;
            3584 : data_o = 1'b0;
            3585 : data_o = 1'b0;
            3586 : data_o = 1'b0;
            3587 : data_o = 1'b0;
            3588 : data_o = 1'b1;
            3589 : data_o = 1'b1;
            3590 : data_o = 1'b1;
            3591 : data_o = 1'b1;
            3592 : data_o = 1'b1;
            3593 : data_o = 1'b1;
            3594 : data_o = 1'b1;
            3595 : data_o = 1'b1;
            3596 : data_o = 1'b1;
            3597 : data_o = 1'b1;
            3598 : data_o = 1'b1;
            3599 : data_o = 1'b1;
            3600 : data_o = 1'b0;
            3601 : data_o = 1'b0;
            3602 : data_o = 1'b0;
            3603 : data_o = 1'b0;
            3604 : data_o = 1'b0;
            3605 : data_o = 1'b0;
            3606 : data_o = 1'b0;
            3607 : data_o = 1'b0;
            3608 : data_o = 1'b0;
            3609 : data_o = 1'b1;
            3610 : data_o = 1'b1;
            3611 : data_o = 1'b1;
            3612 : data_o = 1'b1;
            3613 : data_o = 1'b1;
            3614 : data_o = 1'b1;
            3615 : data_o = 1'b1;
            3616 : data_o = 1'b1;
            3617 : data_o = 1'b1;
            3618 : data_o = 1'b1;
            3619 : data_o = 1'b1;
            3620 : data_o = 1'b1;
            3621 : data_o = 1'b1;
            3622 : data_o = 1'b1;
            3623 : data_o = 1'b0;
            3624 : data_o = 1'b0;
            3625 : data_o = 1'b0;
            3626 : data_o = 1'b0;
            3627 : data_o = 1'b0;
            3628 : data_o = 1'b0;
            3629 : data_o = 1'b0;
            3630 : data_o = 1'b0;
            3631 : data_o = 1'b0;
            3632 : data_o = 1'b1;
            3633 : data_o = 1'b1;
            3634 : data_o = 1'b1;
            3635 : data_o = 1'b1;
            3636 : data_o = 1'b1;
            3637 : data_o = 1'b1;
            3638 : data_o = 1'b1;
            3639 : data_o = 1'b1;
            3640 : data_o = 1'b1;
            3641 : data_o = 1'b1;
            3642 : data_o = 1'b1;
            3643 : data_o = 1'b1;
            3644 : data_o = 1'b1;
            3645 : data_o = 1'b1;
            3646 : data_o = 1'b0;
            3647 : data_o = 1'b0;
            3648 : data_o = 1'b0;
            3649 : data_o = 1'b0;
            3650 : data_o = 1'b0;
            3651 : data_o = 1'b0;
            3652 : data_o = 1'b0;
            3653 : data_o = 1'b1;
            3654 : data_o = 1'b1;
            3655 : data_o = 1'b1;
            3656 : data_o = 1'b1;
            3657 : data_o = 1'b1;
            3658 : data_o = 1'b1;
            3659 : data_o = 1'b1;
            3660 : data_o = 1'b1;
            3661 : data_o = 1'b1;
            3662 : data_o = 1'b1;
            3663 : data_o = 1'b1;
            3664 : data_o = 1'b0;
            3665 : data_o = 1'b0;
            3666 : data_o = 1'b0;
            3667 : data_o = 1'b0;
            3668 : data_o = 1'b0;
            3669 : data_o = 1'b0;
            3670 : data_o = 1'b0;
            3671 : data_o = 1'b0;
            3672 : data_o = 1'b0;
            3673 : data_o = 1'b0;
            3674 : data_o = 1'b0;
            3675 : data_o = 1'b0;
            3676 : data_o = 1'b0;
            3677 : data_o = 1'b0;
            3678 : data_o = 1'b0;
            3679 : data_o = 1'b0;
            3680 : data_o = 1'b0;
            3681 : data_o = 1'b0;
            3682 : data_o = 1'b0;
            3683 : data_o = 1'b0;
            3684 : data_o = 1'b0;
            3685 : data_o = 1'b0;
            3686 : data_o = 1'b0;
            3687 : data_o = 1'b0;
            3688 : data_o = 1'b0;
            3689 : data_o = 1'b0;
            3690 : data_o = 1'b0;
            3691 : data_o = 1'b0;
            3692 : data_o = 1'b0;
            3693 : data_o = 1'b1;
            3694 : data_o = 1'b1;
            3695 : data_o = 1'b1;
            3696 : data_o = 1'b1;
            3697 : data_o = 1'b1;
            3698 : data_o = 1'b1;
            3699 : data_o = 1'b1;
            3700 : data_o = 1'b1;
            3701 : data_o = 1'b1;
            3702 : data_o = 1'b1;
            3703 : data_o = 1'b1;
            3704 : data_o = 1'b1;
            3705 : data_o = 1'b0;
            3706 : data_o = 1'b0;
            3707 : data_o = 1'b0;
            3708 : data_o = 1'b0;
            3709 : data_o = 1'b0;
            3710 : data_o = 1'b0;
            3711 : data_o = 1'b0;
            3712 : data_o = 1'b0;
            3713 : data_o = 1'b0;
            3714 : data_o = 1'b0;
            3715 : data_o = 1'b1;
            3716 : data_o = 1'b1;
            3717 : data_o = 1'b1;
            3718 : data_o = 1'b1;
            3719 : data_o = 1'b1;
            3720 : data_o = 1'b1;
            3721 : data_o = 1'b1;
            3722 : data_o = 1'b1;
            3723 : data_o = 1'b1;
            3724 : data_o = 1'b1;
            3725 : data_o = 1'b1;
            3726 : data_o = 1'b1;
            3727 : data_o = 1'b1;
            3728 : data_o = 1'b0;
            3729 : data_o = 1'b0;
            3730 : data_o = 1'b0;
            3731 : data_o = 1'b0;
            3732 : data_o = 1'b0;
            3733 : data_o = 1'b0;
            3734 : data_o = 1'b0;
            3735 : data_o = 1'b0;
            3736 : data_o = 1'b0;
            3737 : data_o = 1'b0;
            3738 : data_o = 1'b1;
            3739 : data_o = 1'b1;
            3740 : data_o = 1'b1;
            3741 : data_o = 1'b1;
            3742 : data_o = 1'b1;
            3743 : data_o = 1'b1;
            3744 : data_o = 1'b1;
            3745 : data_o = 1'b1;
            3746 : data_o = 1'b1;
            3747 : data_o = 1'b1;
            3748 : data_o = 1'b1;
            3749 : data_o = 1'b1;
            3750 : data_o = 1'b1;
            3751 : data_o = 1'b0;
            3752 : data_o = 1'b0;
            3753 : data_o = 1'b0;
            3754 : data_o = 1'b0;
            3755 : data_o = 1'b0;
            3756 : data_o = 1'b0;
            3757 : data_o = 1'b0;
            3758 : data_o = 1'b0;
            3759 : data_o = 1'b0;
            3760 : data_o = 1'b1;
            3761 : data_o = 1'b1;
            3762 : data_o = 1'b1;
            3763 : data_o = 1'b1;
            3764 : data_o = 1'b1;
            3765 : data_o = 1'b1;
            3766 : data_o = 1'b1;
            3767 : data_o = 1'b1;
            3768 : data_o = 1'b1;
            3769 : data_o = 1'b0;
            3770 : data_o = 1'b0;
            3771 : data_o = 1'b0;
            3772 : data_o = 1'b0;
            3773 : data_o = 1'b0;
            3774 : data_o = 1'b0;
            3775 : data_o = 1'b0;
            3776 : data_o = 1'b0;
            3777 : data_o = 1'b0;
            3778 : data_o = 1'b0;
            3779 : data_o = 1'b0;
            3780 : data_o = 1'b0;
            3781 : data_o = 1'b0;
            3782 : data_o = 1'b0;
            3783 : data_o = 1'b0;
            3784 : data_o = 1'b0;
            3785 : data_o = 1'b0;
            3786 : data_o = 1'b0;
            3787 : data_o = 1'b0;
            3788 : data_o = 1'b0;
            3789 : data_o = 1'b0;
            3790 : data_o = 1'b0;
            3791 : data_o = 1'b0;
            3792 : data_o = 1'b0;
            3793 : data_o = 1'b0;
            3794 : data_o = 1'b0;
            3795 : data_o = 1'b0;
            3796 : data_o = 1'b1;
            3797 : data_o = 1'b1;
            3798 : data_o = 1'b1;
            3799 : data_o = 1'b1;
            3800 : data_o = 1'b1;
            3801 : data_o = 1'b1;
            3802 : data_o = 1'b1;
            3803 : data_o = 1'b1;
            3804 : data_o = 1'b1;
            3805 : data_o = 1'b1;
            3806 : data_o = 1'b1;
            3807 : data_o = 1'b1;
            3808 : data_o = 1'b0;
            3809 : data_o = 1'b0;
            3810 : data_o = 1'b0;
            3811 : data_o = 1'b0;
            3812 : data_o = 1'b0;
            3813 : data_o = 1'b0;
            3814 : data_o = 1'b0;
            3815 : data_o = 1'b0;
            3816 : data_o = 1'b0;
            3817 : data_o = 1'b1;
            3818 : data_o = 1'b1;
            3819 : data_o = 1'b1;
            3820 : data_o = 1'b1;
            3821 : data_o = 1'b1;
            3822 : data_o = 1'b1;
            3823 : data_o = 1'b1;
            3824 : data_o = 1'b1;
            3825 : data_o = 1'b1;
            3826 : data_o = 1'b1;
            3827 : data_o = 1'b1;
            3828 : data_o = 1'b1;
            3829 : data_o = 1'b1;
            3830 : data_o = 1'b1;
            3831 : data_o = 1'b1;
            3832 : data_o = 1'b0;
            3833 : data_o = 1'b0;
            3834 : data_o = 1'b0;
            3835 : data_o = 1'b0;
            3836 : data_o = 1'b0;
            3837 : data_o = 1'b0;
            3838 : data_o = 1'b0;
            3839 : data_o = 1'b0;
            3840 : data_o = 1'b0;
            3841 : data_o = 1'b0;
            3842 : data_o = 1'b1;
            3843 : data_o = 1'b1;
            3844 : data_o = 1'b1;
            3845 : data_o = 1'b1;
            3846 : data_o = 1'b1;
            3847 : data_o = 1'b1;
            3848 : data_o = 1'b1;
            3849 : data_o = 1'b1;
            3850 : data_o = 1'b1;
            3851 : data_o = 1'b1;
            3852 : data_o = 1'b1;
            3853 : data_o = 1'b1;
            3854 : data_o = 1'b1;
            3855 : data_o = 1'b1;
            3856 : data_o = 1'b0;
            3857 : data_o = 1'b0;
            3858 : data_o = 1'b0;
            3859 : data_o = 1'b0;
            3860 : data_o = 1'b0;
            3861 : data_o = 1'b0;
            3862 : data_o = 1'b0;
            3863 : data_o = 1'b0;
            3864 : data_o = 1'b0;
            3865 : data_o = 1'b0;
            3866 : data_o = 1'b0;
            3867 : data_o = 1'b1;
            3868 : data_o = 1'b1;
            3869 : data_o = 1'b1;
            3870 : data_o = 1'b1;
            3871 : data_o = 1'b1;
            3872 : data_o = 1'b1;
            3873 : data_o = 1'b1;
            3874 : data_o = 1'b0;
            3875 : data_o = 1'b0;
            3876 : data_o = 1'b0;
            3877 : data_o = 1'b0;
            3878 : data_o = 1'b0;
            3879 : data_o = 1'b0;
            3880 : data_o = 1'b0;
            3881 : data_o = 1'b0;
            3882 : data_o = 1'b0;
            3883 : data_o = 1'b0;
            3884 : data_o = 1'b0;
            3885 : data_o = 1'b0;
            3886 : data_o = 1'b0;
            3887 : data_o = 1'b0;
            3888 : data_o = 1'b0;
            3889 : data_o = 1'b0;
            3890 : data_o = 1'b0;
            3891 : data_o = 1'b0;
            3892 : data_o = 1'b0;
            3893 : data_o = 1'b0;
            3894 : data_o = 1'b0;
            3895 : data_o = 1'b0;
            3896 : data_o = 1'b0;
            3897 : data_o = 1'b1;
            3898 : data_o = 1'b1;
            3899 : data_o = 1'b1;
            3900 : data_o = 1'b1;
            3901 : data_o = 1'b1;
            3902 : data_o = 1'b1;
            3903 : data_o = 1'b1;
            3904 : data_o = 1'b1;
            3905 : data_o = 1'b1;
            3906 : data_o = 1'b1;
            3907 : data_o = 1'b1;
            3908 : data_o = 1'b1;
            3909 : data_o = 1'b1;
            3910 : data_o = 1'b0;
            3911 : data_o = 1'b0;
            3912 : data_o = 1'b0;
            3913 : data_o = 1'b0;
            3914 : data_o = 1'b0;
            3915 : data_o = 1'b0;
            3916 : data_o = 1'b0;
            3917 : data_o = 1'b0;
            3918 : data_o = 1'b0;
            3919 : data_o = 1'b1;
            3920 : data_o = 1'b1;
            3921 : data_o = 1'b1;
            3922 : data_o = 1'b1;
            3923 : data_o = 1'b1;
            3924 : data_o = 1'b1;
            3925 : data_o = 1'b1;
            3926 : data_o = 1'b1;
            3927 : data_o = 1'b1;
            3928 : data_o = 1'b1;
            3929 : data_o = 1'b1;
            3930 : data_o = 1'b1;
            3931 : data_o = 1'b1;
            3932 : data_o = 1'b1;
            3933 : data_o = 1'b1;
            3934 : data_o = 1'b1;
            3935 : data_o = 1'b0;
            3936 : data_o = 1'b0;
            3937 : data_o = 1'b0;
            3938 : data_o = 1'b0;
            3939 : data_o = 1'b0;
            3940 : data_o = 1'b0;
            3941 : data_o = 1'b0;
            3942 : data_o = 1'b0;
            3943 : data_o = 1'b0;
            3944 : data_o = 1'b0;
            3945 : data_o = 1'b0;
            3946 : data_o = 1'b1;
            3947 : data_o = 1'b1;
            3948 : data_o = 1'b1;
            3949 : data_o = 1'b1;
            3950 : data_o = 1'b1;
            3951 : data_o = 1'b1;
            3952 : data_o = 1'b1;
            3953 : data_o = 1'b1;
            3954 : data_o = 1'b1;
            3955 : data_o = 1'b1;
            3956 : data_o = 1'b1;
            3957 : data_o = 1'b1;
            3958 : data_o = 1'b1;
            3959 : data_o = 1'b1;
            3960 : data_o = 1'b1;
            3961 : data_o = 1'b0;
            3962 : data_o = 1'b0;
            3963 : data_o = 1'b0;
            3964 : data_o = 1'b0;
            3965 : data_o = 1'b0;
            3966 : data_o = 1'b0;
            3967 : data_o = 1'b0;
            3968 : data_o = 1'b0;
            3969 : data_o = 1'b0;
            3970 : data_o = 1'b0;
            3971 : data_o = 1'b0;
            3972 : data_o = 1'b0;
            3973 : data_o = 1'b0;
            3974 : data_o = 1'b1;
            3975 : data_o = 1'b1;
            3976 : data_o = 1'b1;
            3977 : data_o = 1'b0;
            3978 : data_o = 1'b0;
            3979 : data_o = 1'b0;
            3980 : data_o = 1'b0;
            3981 : data_o = 1'b0;
            3982 : data_o = 1'b0;
            3983 : data_o = 1'b0;
            3984 : data_o = 1'b0;
            3985 : data_o = 1'b0;
            3986 : data_o = 1'b0;
            3987 : data_o = 1'b0;
            3988 : data_o = 1'b0;
            3989 : data_o = 1'b0;
            3990 : data_o = 1'b0;
            3991 : data_o = 1'b0;
            3992 : data_o = 1'b0;
            3993 : data_o = 1'b0;
            3994 : data_o = 1'b0;
            3995 : data_o = 1'b0;
            3996 : data_o = 1'b0;
            3997 : data_o = 1'b0;
            3998 : data_o = 1'b0;
            3999 : data_o = 1'b1;
            4000 : data_o = 1'b1;
            4001 : data_o = 1'b1;
            4002 : data_o = 1'b1;
            4003 : data_o = 1'b1;
            4004 : data_o = 1'b1;
            4005 : data_o = 1'b1;
            4006 : data_o = 1'b1;
            4007 : data_o = 1'b1;
            4008 : data_o = 1'b1;
            4009 : data_o = 1'b1;
            4010 : data_o = 1'b1;
            4011 : data_o = 1'b1;
            4012 : data_o = 1'b0;
            4013 : data_o = 1'b0;
            4014 : data_o = 1'b0;
            4015 : data_o = 1'b0;
            4016 : data_o = 1'b0;
            4017 : data_o = 1'b0;
            4018 : data_o = 1'b0;
            4019 : data_o = 1'b0;
            4020 : data_o = 1'b0;
            4021 : data_o = 1'b1;
            4022 : data_o = 1'b1;
            4023 : data_o = 1'b1;
            4024 : data_o = 1'b1;
            4025 : data_o = 1'b1;
            4026 : data_o = 1'b1;
            4027 : data_o = 1'b1;
            4028 : data_o = 1'b1;
            4029 : data_o = 1'b1;
            4030 : data_o = 1'b1;
            4031 : data_o = 1'b1;
            4032 : data_o = 1'b1;
            4033 : data_o = 1'b1;
            4034 : data_o = 1'b1;
            4035 : data_o = 1'b1;
            4036 : data_o = 1'b1;
            4037 : data_o = 1'b1;
            4038 : data_o = 1'b1;
            4039 : data_o = 1'b0;
            4040 : data_o = 1'b0;
            4041 : data_o = 1'b0;
            4042 : data_o = 1'b0;
            4043 : data_o = 1'b0;
            4044 : data_o = 1'b0;
            4045 : data_o = 1'b0;
            4046 : data_o = 1'b0;
            4047 : data_o = 1'b0;
            4048 : data_o = 1'b0;
            4049 : data_o = 1'b1;
            4050 : data_o = 1'b1;
            4051 : data_o = 1'b1;
            4052 : data_o = 1'b1;
            4053 : data_o = 1'b1;
            4054 : data_o = 1'b1;
            4055 : data_o = 1'b1;
            4056 : data_o = 1'b1;
            4057 : data_o = 1'b1;
            4058 : data_o = 1'b1;
            4059 : data_o = 1'b1;
            4060 : data_o = 1'b1;
            4061 : data_o = 1'b1;
            4062 : data_o = 1'b1;
            4063 : data_o = 1'b1;
            4064 : data_o = 1'b1;
            4065 : data_o = 1'b0;
            4066 : data_o = 1'b0;
            4067 : data_o = 1'b0;
            4068 : data_o = 1'b0;
            4069 : data_o = 1'b0;
            4070 : data_o = 1'b0;
            4071 : data_o = 1'b0;
            4072 : data_o = 1'b0;
            4073 : data_o = 1'b0;
            4074 : data_o = 1'b0;
            4075 : data_o = 1'b0;
            4076 : data_o = 1'b0;
            4077 : data_o = 1'b0;
            4078 : data_o = 1'b0;
            4079 : data_o = 1'b0;
            4080 : data_o = 1'b0;
            4081 : data_o = 1'b0;
            4082 : data_o = 1'b0;
            4083 : data_o = 1'b0;
            4084 : data_o = 1'b0;
            4085 : data_o = 1'b0;
            4086 : data_o = 1'b0;
            4087 : data_o = 1'b0;
            4088 : data_o = 1'b0;
            4089 : data_o = 1'b0;
            4090 : data_o = 1'b0;
            4091 : data_o = 1'b0;
            4092 : data_o = 1'b0;
            4093 : data_o = 1'b0;
            4094 : data_o = 1'b0;
            4095 : data_o = 1'b0;
            4096 : data_o = 1'b0;
            4097 : data_o = 1'b0;
            4098 : data_o = 1'b0;
            4099 : data_o = 1'b0;
            4100 : data_o = 1'b1;
            4101 : data_o = 1'b1;
            4102 : data_o = 1'b1;
            4103 : data_o = 1'b1;
            4104 : data_o = 1'b1;
            4105 : data_o = 1'b1;
            4106 : data_o = 1'b1;
            4107 : data_o = 1'b1;
            4108 : data_o = 1'b1;
            4109 : data_o = 1'b1;
            4110 : data_o = 1'b1;
            4111 : data_o = 1'b1;
            4112 : data_o = 1'b1;
            4113 : data_o = 1'b1;
            4114 : data_o = 1'b1;
            4115 : data_o = 1'b0;
            4116 : data_o = 1'b0;
            4117 : data_o = 1'b0;
            4118 : data_o = 1'b0;
            4119 : data_o = 1'b0;
            4120 : data_o = 1'b0;
            4121 : data_o = 1'b0;
            4122 : data_o = 1'b0;
            4123 : data_o = 1'b1;
            4124 : data_o = 1'b1;
            4125 : data_o = 1'b1;
            4126 : data_o = 1'b1;
            4127 : data_o = 1'b1;
            4128 : data_o = 1'b1;
            4129 : data_o = 1'b1;
            4130 : data_o = 1'b1;
            4131 : data_o = 1'b1;
            4132 : data_o = 1'b1;
            4133 : data_o = 1'b1;
            4134 : data_o = 1'b1;
            4135 : data_o = 1'b1;
            4136 : data_o = 1'b1;
            4137 : data_o = 1'b1;
            4138 : data_o = 1'b1;
            4139 : data_o = 1'b1;
            4140 : data_o = 1'b1;
            4141 : data_o = 1'b1;
            4142 : data_o = 1'b1;
            4143 : data_o = 1'b1;
            4144 : data_o = 1'b1;
            4145 : data_o = 1'b1;
            4146 : data_o = 1'b1;
            4147 : data_o = 1'b1;
            4148 : data_o = 1'b0;
            4149 : data_o = 1'b0;
            4150 : data_o = 1'b0;
            4151 : data_o = 1'b1;
            4152 : data_o = 1'b1;
            4153 : data_o = 1'b1;
            4154 : data_o = 1'b1;
            4155 : data_o = 1'b1;
            4156 : data_o = 1'b1;
            4157 : data_o = 1'b1;
            4158 : data_o = 1'b1;
            4159 : data_o = 1'b1;
            4160 : data_o = 1'b1;
            4161 : data_o = 1'b1;
            4162 : data_o = 1'b1;
            4163 : data_o = 1'b1;
            4164 : data_o = 1'b1;
            4165 : data_o = 1'b1;
            4166 : data_o = 1'b1;
            4167 : data_o = 1'b1;
            4168 : data_o = 1'b1;
            4169 : data_o = 1'b0;
            4170 : data_o = 1'b0;
            4171 : data_o = 1'b0;
            4172 : data_o = 1'b0;
            4173 : data_o = 1'b0;
            4174 : data_o = 1'b0;
            4175 : data_o = 1'b0;
            4176 : data_o = 1'b0;
            4177 : data_o = 1'b0;
            4178 : data_o = 1'b0;
            4179 : data_o = 1'b0;
            4180 : data_o = 1'b0;
            4181 : data_o = 1'b0;
            4182 : data_o = 1'b0;
            4183 : data_o = 1'b0;
            4184 : data_o = 1'b0;
            4185 : data_o = 1'b0;
            4186 : data_o = 1'b0;
            4187 : data_o = 1'b0;
            4188 : data_o = 1'b0;
            4189 : data_o = 1'b0;
            4190 : data_o = 1'b0;
            4191 : data_o = 1'b0;
            4192 : data_o = 1'b0;
            4193 : data_o = 1'b0;
            4194 : data_o = 1'b0;
            4195 : data_o = 1'b0;
            4196 : data_o = 1'b0;
            4197 : data_o = 1'b0;
            4198 : data_o = 1'b0;
            4199 : data_o = 1'b0;
            4200 : data_o = 1'b0;
            4201 : data_o = 1'b0;
            4202 : data_o = 1'b0;
            4203 : data_o = 1'b1;
            4204 : data_o = 1'b1;
            4205 : data_o = 1'b1;
            4206 : data_o = 1'b1;
            4207 : data_o = 1'b1;
            4208 : data_o = 1'b1;
            4209 : data_o = 1'b1;
            4210 : data_o = 1'b1;
            4211 : data_o = 1'b1;
            4212 : data_o = 1'b1;
            4213 : data_o = 1'b1;
            4214 : data_o = 1'b1;
            4215 : data_o = 1'b1;
            4216 : data_o = 1'b1;
            4217 : data_o = 1'b1;
            4218 : data_o = 1'b1;
            4219 : data_o = 1'b1;
            4220 : data_o = 1'b1;
            4221 : data_o = 1'b1;
            4222 : data_o = 1'b1;
            4223 : data_o = 1'b1;
            4224 : data_o = 1'b1;
            4225 : data_o = 1'b1;
            4226 : data_o = 1'b1;
            4227 : data_o = 1'b1;
            4228 : data_o = 1'b1;
            4229 : data_o = 1'b1;
            4230 : data_o = 1'b1;
            4231 : data_o = 1'b1;
            4232 : data_o = 1'b1;
            4233 : data_o = 1'b1;
            4234 : data_o = 1'b1;
            4235 : data_o = 1'b1;
            4236 : data_o = 1'b1;
            4237 : data_o = 1'b1;
            4238 : data_o = 1'b1;
            4239 : data_o = 1'b1;
            4240 : data_o = 1'b1;
            4241 : data_o = 1'b1;
            4242 : data_o = 1'b1;
            4243 : data_o = 1'b1;
            4244 : data_o = 1'b1;
            4245 : data_o = 1'b1;
            4246 : data_o = 1'b1;
            4247 : data_o = 1'b1;
            4248 : data_o = 1'b1;
            4249 : data_o = 1'b1;
            4250 : data_o = 1'b1;
            4251 : data_o = 1'b1;
            4252 : data_o = 1'b1;
            4253 : data_o = 1'b1;
            4254 : data_o = 1'b0;
            4255 : data_o = 1'b0;
            4256 : data_o = 1'b0;
            4257 : data_o = 1'b1;
            4258 : data_o = 1'b1;
            4259 : data_o = 1'b1;
            4260 : data_o = 1'b1;
            4261 : data_o = 1'b1;
            4262 : data_o = 1'b1;
            4263 : data_o = 1'b1;
            4264 : data_o = 1'b1;
            4265 : data_o = 1'b1;
            4266 : data_o = 1'b1;
            4267 : data_o = 1'b1;
            4268 : data_o = 1'b1;
            4269 : data_o = 1'b1;
            4270 : data_o = 1'b1;
            4271 : data_o = 1'b1;
            4272 : data_o = 1'b1;
            4273 : data_o = 1'b1;
            4274 : data_o = 1'b0;
            4275 : data_o = 1'b0;
            4276 : data_o = 1'b0;
            4277 : data_o = 1'b0;
            4278 : data_o = 1'b0;
            4279 : data_o = 1'b0;
            4280 : data_o = 1'b0;
            4281 : data_o = 1'b0;
            4282 : data_o = 1'b0;
            4283 : data_o = 1'b0;
            4284 : data_o = 1'b0;
            4285 : data_o = 1'b0;
            4286 : data_o = 1'b0;
            4287 : data_o = 1'b0;
            4288 : data_o = 1'b0;
            4289 : data_o = 1'b0;
            4290 : data_o = 1'b0;
            4291 : data_o = 1'b0;
            4292 : data_o = 1'b0;
            4293 : data_o = 1'b0;
            4294 : data_o = 1'b0;
            4295 : data_o = 1'b0;
            4296 : data_o = 1'b0;
            4297 : data_o = 1'b0;
            4298 : data_o = 1'b0;
            4299 : data_o = 1'b0;
            4300 : data_o = 1'b0;
            4301 : data_o = 1'b0;
            4302 : data_o = 1'b0;
            4303 : data_o = 1'b0;
            4304 : data_o = 1'b0;
            4305 : data_o = 1'b0;
            4306 : data_o = 1'b1;
            4307 : data_o = 1'b1;
            4308 : data_o = 1'b1;
            4309 : data_o = 1'b1;
            4310 : data_o = 1'b1;
            4311 : data_o = 1'b1;
            4312 : data_o = 1'b1;
            4313 : data_o = 1'b1;
            4314 : data_o = 1'b1;
            4315 : data_o = 1'b1;
            4316 : data_o = 1'b1;
            4317 : data_o = 1'b1;
            4318 : data_o = 1'b1;
            4319 : data_o = 1'b1;
            4320 : data_o = 1'b1;
            4321 : data_o = 1'b1;
            4322 : data_o = 1'b1;
            4323 : data_o = 1'b1;
            4324 : data_o = 1'b1;
            4325 : data_o = 1'b1;
            4326 : data_o = 1'b1;
            4327 : data_o = 1'b1;
            4328 : data_o = 1'b1;
            4329 : data_o = 1'b1;
            4330 : data_o = 1'b1;
            4331 : data_o = 1'b1;
            4332 : data_o = 1'b1;
            4333 : data_o = 1'b1;
            4334 : data_o = 1'b1;
            4335 : data_o = 1'b1;
            4336 : data_o = 1'b1;
            4337 : data_o = 1'b1;
            4338 : data_o = 1'b1;
            4339 : data_o = 1'b1;
            4340 : data_o = 1'b1;
            4341 : data_o = 1'b1;
            4342 : data_o = 1'b1;
            4343 : data_o = 1'b1;
            4344 : data_o = 1'b1;
            4345 : data_o = 1'b1;
            4346 : data_o = 1'b1;
            4347 : data_o = 1'b1;
            4348 : data_o = 1'b1;
            4349 : data_o = 1'b1;
            4350 : data_o = 1'b1;
            4351 : data_o = 1'b1;
            4352 : data_o = 1'b1;
            4353 : data_o = 1'b1;
            4354 : data_o = 1'b1;
            4355 : data_o = 1'b1;
            4356 : data_o = 1'b1;
            4357 : data_o = 1'b1;
            4358 : data_o = 1'b1;
            4359 : data_o = 1'b1;
            4360 : data_o = 1'b1;
            4361 : data_o = 1'b1;
            4362 : data_o = 1'b1;
            4363 : data_o = 1'b1;
            4364 : data_o = 1'b1;
            4365 : data_o = 1'b1;
            4366 : data_o = 1'b1;
            4367 : data_o = 1'b1;
            4368 : data_o = 1'b1;
            4369 : data_o = 1'b1;
            4370 : data_o = 1'b1;
            4371 : data_o = 1'b1;
            4372 : data_o = 1'b1;
            4373 : data_o = 1'b1;
            4374 : data_o = 1'b1;
            4375 : data_o = 1'b1;
            4376 : data_o = 1'b1;
            4377 : data_o = 1'b0;
            4378 : data_o = 1'b0;
            4379 : data_o = 1'b0;
            4380 : data_o = 1'b0;
            4381 : data_o = 1'b0;
            4382 : data_o = 1'b0;
            4383 : data_o = 1'b0;
            4384 : data_o = 1'b0;
            4385 : data_o = 1'b0;
            4386 : data_o = 1'b0;
            4387 : data_o = 1'b0;
            4388 : data_o = 1'b0;
            4389 : data_o = 1'b0;
            4390 : data_o = 1'b0;
            4391 : data_o = 1'b0;
            4392 : data_o = 1'b0;
            4393 : data_o = 1'b0;
            4394 : data_o = 1'b0;
            4395 : data_o = 1'b0;
            4396 : data_o = 1'b0;
            4397 : data_o = 1'b0;
            4398 : data_o = 1'b0;
            4399 : data_o = 1'b0;
            4400 : data_o = 1'b0;
            4401 : data_o = 1'b0;
            4402 : data_o = 1'b0;
            4403 : data_o = 1'b0;
            4404 : data_o = 1'b0;
            4405 : data_o = 1'b0;
            4406 : data_o = 1'b0;
            4407 : data_o = 1'b0;
            4408 : data_o = 1'b0;
            4409 : data_o = 1'b0;
            4410 : data_o = 1'b0;
            4411 : data_o = 1'b1;
            4412 : data_o = 1'b1;
            4413 : data_o = 1'b1;
            4414 : data_o = 1'b1;
            4415 : data_o = 1'b1;
            4416 : data_o = 1'b1;
            4417 : data_o = 1'b1;
            4418 : data_o = 1'b0;
            4419 : data_o = 1'b0;
            4420 : data_o = 1'b0;
            4421 : data_o = 1'b0;
            4422 : data_o = 1'b0;
            4423 : data_o = 1'b0;
            4424 : data_o = 1'b1;
            4425 : data_o = 1'b1;
            4426 : data_o = 1'b1;
            4427 : data_o = 1'b1;
            4428 : data_o = 1'b1;
            4429 : data_o = 1'b1;
            4430 : data_o = 1'b1;
            4431 : data_o = 1'b1;
            4432 : data_o = 1'b1;
            4433 : data_o = 1'b1;
            4434 : data_o = 1'b1;
            4435 : data_o = 1'b1;
            4436 : data_o = 1'b1;
            4437 : data_o = 1'b1;
            4438 : data_o = 1'b1;
            4439 : data_o = 1'b1;
            4440 : data_o = 1'b1;
            4441 : data_o = 1'b1;
            4442 : data_o = 1'b1;
            4443 : data_o = 1'b1;
            4444 : data_o = 1'b1;
            4445 : data_o = 1'b1;
            4446 : data_o = 1'b1;
            4447 : data_o = 1'b1;
            4448 : data_o = 1'b1;
            4449 : data_o = 1'b1;
            4450 : data_o = 1'b1;
            4451 : data_o = 1'b1;
            4452 : data_o = 1'b1;
            4453 : data_o = 1'b1;
            4454 : data_o = 1'b1;
            4455 : data_o = 1'b1;
            4456 : data_o = 1'b1;
            4457 : data_o = 1'b1;
            4458 : data_o = 1'b1;
            4459 : data_o = 1'b1;
            4460 : data_o = 1'b1;
            4461 : data_o = 1'b1;
            4462 : data_o = 1'b1;
            4463 : data_o = 1'b1;
            4464 : data_o = 1'b1;
            4465 : data_o = 1'b1;
            4466 : data_o = 1'b1;
            4467 : data_o = 1'b1;
            4468 : data_o = 1'b1;
            4469 : data_o = 1'b1;
            4470 : data_o = 1'b1;
            4471 : data_o = 1'b1;
            4472 : data_o = 1'b1;
            4473 : data_o = 1'b1;
            4474 : data_o = 1'b1;
            4475 : data_o = 1'b1;
            4476 : data_o = 1'b1;
            4477 : data_o = 1'b1;
            4478 : data_o = 1'b1;
            4479 : data_o = 1'b1;
            4480 : data_o = 1'b0;
            4481 : data_o = 1'b0;
            4482 : data_o = 1'b0;
            4483 : data_o = 1'b0;
            4484 : data_o = 1'b0;
            4485 : data_o = 1'b0;
            4486 : data_o = 1'b0;
            4487 : data_o = 1'b0;
            4488 : data_o = 1'b0;
            4489 : data_o = 1'b0;
            4490 : data_o = 1'b0;
            4491 : data_o = 1'b0;
            4492 : data_o = 1'b0;
            4493 : data_o = 1'b0;
            4494 : data_o = 1'b0;
            4495 : data_o = 1'b0;
            4496 : data_o = 1'b0;
            4497 : data_o = 1'b0;
            4498 : data_o = 1'b0;
            4499 : data_o = 1'b0;
            4500 : data_o = 1'b0;
            4501 : data_o = 1'b0;
            4502 : data_o = 1'b0;
            4503 : data_o = 1'b0;
            4504 : data_o = 1'b0;
            4505 : data_o = 1'b0;
            4506 : data_o = 1'b0;
            4507 : data_o = 1'b0;
            4508 : data_o = 1'b0;
            4509 : data_o = 1'b0;
            4510 : data_o = 1'b0;
            4511 : data_o = 1'b0;
            4512 : data_o = 1'b0;
            4513 : data_o = 1'b0;
            4514 : data_o = 1'b0;
            4515 : data_o = 1'b0;
            4516 : data_o = 1'b1;
            4517 : data_o = 1'b1;
            4518 : data_o = 1'b1;
            4519 : data_o = 1'b1;
            4520 : data_o = 1'b1;
            4521 : data_o = 1'b0;
            4522 : data_o = 1'b0;
            4523 : data_o = 1'b0;
            4524 : data_o = 1'b0;
            4525 : data_o = 1'b0;
            4526 : data_o = 1'b0;
            4527 : data_o = 1'b0;
            4528 : data_o = 1'b0;
            4529 : data_o = 1'b1;
            4530 : data_o = 1'b1;
            4531 : data_o = 1'b1;
            4532 : data_o = 1'b1;
            4533 : data_o = 1'b1;
            4534 : data_o = 1'b1;
            4535 : data_o = 1'b1;
            4536 : data_o = 1'b1;
            4537 : data_o = 1'b1;
            4538 : data_o = 1'b1;
            4539 : data_o = 1'b1;
            4540 : data_o = 1'b1;
            4541 : data_o = 1'b1;
            4542 : data_o = 1'b1;
            4543 : data_o = 1'b1;
            4544 : data_o = 1'b1;
            4545 : data_o = 1'b1;
            4546 : data_o = 1'b1;
            4547 : data_o = 1'b1;
            4548 : data_o = 1'b1;
            4549 : data_o = 1'b1;
            4550 : data_o = 1'b1;
            4551 : data_o = 1'b1;
            4552 : data_o = 1'b1;
            4553 : data_o = 1'b1;
            4554 : data_o = 1'b1;
            4555 : data_o = 1'b1;
            4556 : data_o = 1'b1;
            4557 : data_o = 1'b1;
            4558 : data_o = 1'b1;
            4559 : data_o = 1'b1;
            4560 : data_o = 1'b1;
            4561 : data_o = 1'b1;
            4562 : data_o = 1'b1;
            4563 : data_o = 1'b1;
            4564 : data_o = 1'b1;
            4565 : data_o = 1'b1;
            4566 : data_o = 1'b1;
            4567 : data_o = 1'b1;
            4568 : data_o = 1'b1;
            4569 : data_o = 1'b1;
            4570 : data_o = 1'b1;
            4571 : data_o = 1'b1;
            4572 : data_o = 1'b1;
            4573 : data_o = 1'b1;
            4574 : data_o = 1'b1;
            4575 : data_o = 1'b1;
            4576 : data_o = 1'b1;
            4577 : data_o = 1'b1;
            4578 : data_o = 1'b1;
            4579 : data_o = 1'b1;
            4580 : data_o = 1'b1;
            4581 : data_o = 1'b1;
            4582 : data_o = 1'b1;
            4583 : data_o = 1'b1;
            4584 : data_o = 1'b0;
            4585 : data_o = 1'b0;
            4586 : data_o = 1'b0;
            4587 : data_o = 1'b0;
            4588 : data_o = 1'b0;
            4589 : data_o = 1'b0;
            4590 : data_o = 1'b0;
            4591 : data_o = 1'b0;
            4592 : data_o = 1'b0;
            4593 : data_o = 1'b0;
            4594 : data_o = 1'b0;
            4595 : data_o = 1'b0;
            4596 : data_o = 1'b0;
            4597 : data_o = 1'b0;
            4598 : data_o = 1'b0;
            4599 : data_o = 1'b0;
            4600 : data_o = 1'b0;
            4601 : data_o = 1'b0;
            4602 : data_o = 1'b0;
            4603 : data_o = 1'b0;
            4604 : data_o = 1'b0;
            4605 : data_o = 1'b0;
            4606 : data_o = 1'b0;
            4607 : data_o = 1'b0;
            4608 : data_o = 1'b0;
            4609 : data_o = 1'b0;
            4610 : data_o = 1'b0;
            4611 : data_o = 1'b0;
            4612 : data_o = 1'b0;
            4613 : data_o = 1'b0;
            4614 : data_o = 1'b0;
            4615 : data_o = 1'b0;
            4616 : data_o = 1'b0;
            4617 : data_o = 1'b0;
            4618 : data_o = 1'b0;
            4619 : data_o = 1'b0;
            4620 : data_o = 1'b0;
            4621 : data_o = 1'b0;
            4622 : data_o = 1'b1;
            4623 : data_o = 1'b1;
            4624 : data_o = 1'b1;
            4625 : data_o = 1'b0;
            4626 : data_o = 1'b0;
            4627 : data_o = 1'b0;
            4628 : data_o = 1'b0;
            4629 : data_o = 1'b0;
            4630 : data_o = 1'b0;
            4631 : data_o = 1'b0;
            4632 : data_o = 1'b0;
            4633 : data_o = 1'b0;
            4634 : data_o = 1'b0;
            4635 : data_o = 1'b1;
            4636 : data_o = 1'b1;
            4637 : data_o = 1'b1;
            4638 : data_o = 1'b1;
            4639 : data_o = 1'b1;
            4640 : data_o = 1'b1;
            4641 : data_o = 1'b1;
            4642 : data_o = 1'b1;
            4643 : data_o = 1'b1;
            4644 : data_o = 1'b1;
            4645 : data_o = 1'b1;
            4646 : data_o = 1'b1;
            4647 : data_o = 1'b1;
            4648 : data_o = 1'b1;
            4649 : data_o = 1'b1;
            4650 : data_o = 1'b1;
            4651 : data_o = 1'b1;
            4652 : data_o = 1'b1;
            4653 : data_o = 1'b1;
            4654 : data_o = 1'b1;
            4655 : data_o = 1'b1;
            4656 : data_o = 1'b1;
            4657 : data_o = 1'b1;
            4658 : data_o = 1'b1;
            4659 : data_o = 1'b1;
            4660 : data_o = 1'b1;
            4661 : data_o = 1'b1;
            4662 : data_o = 1'b1;
            4663 : data_o = 1'b1;
            4664 : data_o = 1'b1;
            4665 : data_o = 1'b1;
            4666 : data_o = 1'b1;
            4667 : data_o = 1'b1;
            4668 : data_o = 1'b1;
            4669 : data_o = 1'b1;
            4670 : data_o = 1'b1;
            4671 : data_o = 1'b1;
            4672 : data_o = 1'b1;
            4673 : data_o = 1'b1;
            4674 : data_o = 1'b1;
            4675 : data_o = 1'b1;
            4676 : data_o = 1'b1;
            4677 : data_o = 1'b1;
            4678 : data_o = 1'b1;
            4679 : data_o = 1'b1;
            4680 : data_o = 1'b1;
            4681 : data_o = 1'b1;
            4682 : data_o = 1'b1;
            4683 : data_o = 1'b1;
            4684 : data_o = 1'b1;
            4685 : data_o = 1'b1;
            4686 : data_o = 1'b1;
            4687 : data_o = 1'b1;
            4688 : data_o = 1'b0;
            4689 : data_o = 1'b0;
            4690 : data_o = 1'b0;
            4691 : data_o = 1'b0;
            4692 : data_o = 1'b0;
            4693 : data_o = 1'b0;
            4694 : data_o = 1'b0;
            4695 : data_o = 1'b0;
            4696 : data_o = 1'b0;
            4697 : data_o = 1'b0;
            4698 : data_o = 1'b0;
            4699 : data_o = 1'b0;
            4700 : data_o = 1'b0;
            4701 : data_o = 1'b0;
            4702 : data_o = 1'b0;
            4703 : data_o = 1'b0;
            4704 : data_o = 1'b0;
            4705 : data_o = 1'b0;
            4706 : data_o = 1'b0;
            4707 : data_o = 1'b0;
            4708 : data_o = 1'b0;
            4709 : data_o = 1'b0;
            4710 : data_o = 1'b0;
            4711 : data_o = 1'b0;
            4712 : data_o = 1'b0;
            4713 : data_o = 1'b0;
            4714 : data_o = 1'b0;
            4715 : data_o = 1'b0;
            4716 : data_o = 1'b0;
            4717 : data_o = 1'b0;
            4718 : data_o = 1'b0;
            4719 : data_o = 1'b0;
            4720 : data_o = 1'b0;
            4721 : data_o = 1'b0;
            4722 : data_o = 1'b0;
            4723 : data_o = 1'b0;
            4724 : data_o = 1'b0;
            4725 : data_o = 1'b0;
            4726 : data_o = 1'b1;
            4727 : data_o = 1'b1;
            4728 : data_o = 1'b1;
            4729 : data_o = 1'b0;
            4730 : data_o = 1'b0;
            4731 : data_o = 1'b0;
            4732 : data_o = 1'b0;
            4733 : data_o = 1'b0;
            4734 : data_o = 1'b0;
            4735 : data_o = 1'b0;
            4736 : data_o = 1'b0;
            4737 : data_o = 1'b0;
            4738 : data_o = 1'b0;
            4739 : data_o = 1'b0;
            4740 : data_o = 1'b1;
            4741 : data_o = 1'b1;
            4742 : data_o = 1'b1;
            4743 : data_o = 1'b1;
            4744 : data_o = 1'b1;
            4745 : data_o = 1'b1;
            4746 : data_o = 1'b1;
            4747 : data_o = 1'b1;
            4748 : data_o = 1'b1;
            4749 : data_o = 1'b1;
            4750 : data_o = 1'b1;
            4751 : data_o = 1'b1;
            4752 : data_o = 1'b1;
            4753 : data_o = 1'b1;
            4754 : data_o = 1'b1;
            4755 : data_o = 1'b1;
            4756 : data_o = 1'b1;
            4757 : data_o = 1'b1;
            4758 : data_o = 1'b1;
            4759 : data_o = 1'b1;
            4760 : data_o = 1'b1;
            4761 : data_o = 1'b1;
            4762 : data_o = 1'b1;
            4763 : data_o = 1'b1;
            4764 : data_o = 1'b1;
            4765 : data_o = 1'b1;
            4766 : data_o = 1'b1;
            4767 : data_o = 1'b1;
            4768 : data_o = 1'b1;
            4769 : data_o = 1'b1;
            4770 : data_o = 1'b1;
            4771 : data_o = 1'b1;
            4772 : data_o = 1'b1;
            4773 : data_o = 1'b1;
            4774 : data_o = 1'b1;
            4775 : data_o = 1'b1;
            4776 : data_o = 1'b1;
            4777 : data_o = 1'b1;
            4778 : data_o = 1'b1;
            4779 : data_o = 1'b1;
            4780 : data_o = 1'b1;
            4781 : data_o = 1'b1;
            4782 : data_o = 1'b1;
            4783 : data_o = 1'b1;
            4784 : data_o = 1'b1;
            4785 : data_o = 1'b1;
            4786 : data_o = 1'b1;
            4787 : data_o = 1'b1;
            4788 : data_o = 1'b1;
            4789 : data_o = 1'b1;
            4790 : data_o = 1'b1;
            4791 : data_o = 1'b1;
            4792 : data_o = 1'b1;
            4793 : data_o = 1'b0;
            4794 : data_o = 1'b0;
            4795 : data_o = 1'b0;
            4796 : data_o = 1'b0;
            4797 : data_o = 1'b0;
            4798 : data_o = 1'b0;
            4799 : data_o = 1'b0;
            4800 : data_o = 1'b0;
            4801 : data_o = 1'b0;
            4802 : data_o = 1'b0;
            4803 : data_o = 1'b0;
            4804 : data_o = 1'b0;
            4805 : data_o = 1'b0;
            4806 : data_o = 1'b0;
            4807 : data_o = 1'b0;
            4808 : data_o = 1'b0;
            4809 : data_o = 1'b0;
            4810 : data_o = 1'b0;
            4811 : data_o = 1'b0;
            4812 : data_o = 1'b0;
            4813 : data_o = 1'b0;
            4814 : data_o = 1'b0;
            4815 : data_o = 1'b0;
            4816 : data_o = 1'b0;
            4817 : data_o = 1'b0;
            4818 : data_o = 1'b0;
            4819 : data_o = 1'b0;
            4820 : data_o = 1'b0;
            4821 : data_o = 1'b0;
            4822 : data_o = 1'b0;
            4823 : data_o = 1'b0;
            4824 : data_o = 1'b0;
            4825 : data_o = 1'b0;
            4826 : data_o = 1'b0;
            4827 : data_o = 1'b0;
            4828 : data_o = 1'b0;
            4829 : data_o = 1'b0;
            4830 : data_o = 1'b0;
            4831 : data_o = 1'b0;
            4832 : data_o = 1'b0;
            4833 : data_o = 1'b0;
            4834 : data_o = 1'b0;
            4835 : data_o = 1'b0;
            4836 : data_o = 1'b0;
            4837 : data_o = 1'b0;
            4838 : data_o = 1'b0;
            4839 : data_o = 1'b0;
            4840 : data_o = 1'b0;
            4841 : data_o = 1'b0;
            4842 : data_o = 1'b0;
            4843 : data_o = 1'b0;
            4844 : data_o = 1'b0;
            4845 : data_o = 1'b0;
            4846 : data_o = 1'b1;
            4847 : data_o = 1'b1;
            4848 : data_o = 1'b1;
            4849 : data_o = 1'b1;
            4850 : data_o = 1'b1;
            4851 : data_o = 1'b1;
            4852 : data_o = 1'b1;
            4853 : data_o = 1'b1;
            4854 : data_o = 1'b1;
            4855 : data_o = 1'b1;
            4856 : data_o = 1'b1;
            4857 : data_o = 1'b1;
            4858 : data_o = 1'b1;
            4859 : data_o = 1'b1;
            4860 : data_o = 1'b1;
            4861 : data_o = 1'b1;
            4862 : data_o = 1'b1;
            4863 : data_o = 1'b1;
            4864 : data_o = 1'b1;
            4865 : data_o = 1'b1;
            4866 : data_o = 1'b1;
            4867 : data_o = 1'b1;
            4868 : data_o = 1'b1;
            4869 : data_o = 1'b1;
            4870 : data_o = 1'b1;
            4871 : data_o = 1'b1;
            4872 : data_o = 1'b1;
            4873 : data_o = 1'b1;
            4874 : data_o = 1'b1;
            4875 : data_o = 1'b1;
            4876 : data_o = 1'b1;
            4877 : data_o = 1'b1;
            4878 : data_o = 1'b1;
            4879 : data_o = 1'b1;
            4880 : data_o = 1'b1;
            4881 : data_o = 1'b1;
            4882 : data_o = 1'b1;
            4883 : data_o = 1'b1;
            4884 : data_o = 1'b1;
            4885 : data_o = 1'b1;
            4886 : data_o = 1'b1;
            4887 : data_o = 1'b1;
            4888 : data_o = 1'b1;
            4889 : data_o = 1'b1;
            4890 : data_o = 1'b1;
            4891 : data_o = 1'b1;
            4892 : data_o = 1'b1;
            4893 : data_o = 1'b1;
            4894 : data_o = 1'b1;
            4895 : data_o = 1'b1;
            4896 : data_o = 1'b1;
            4897 : data_o = 1'b1;
            4898 : data_o = 1'b0;
            4899 : data_o = 1'b0;
            4900 : data_o = 1'b0;
            4901 : data_o = 1'b0;
            4902 : data_o = 1'b0;
            4903 : data_o = 1'b0;
            4904 : data_o = 1'b0;
            4905 : data_o = 1'b0;
            4906 : data_o = 1'b0;
            4907 : data_o = 1'b0;
            4908 : data_o = 1'b0;
            4909 : data_o = 1'b0;
            4910 : data_o = 1'b0;
            4911 : data_o = 1'b0;
            4912 : data_o = 1'b0;
            4913 : data_o = 1'b0;
            4914 : data_o = 1'b0;
            4915 : data_o = 1'b0;
            4916 : data_o = 1'b0;
            4917 : data_o = 1'b0;
            4918 : data_o = 1'b0;
            4919 : data_o = 1'b0;
            4920 : data_o = 1'b0;
            4921 : data_o = 1'b0;
            4922 : data_o = 1'b0;
            4923 : data_o = 1'b0;
            4924 : data_o = 1'b0;
            4925 : data_o = 1'b0;
            4926 : data_o = 1'b0;
            4927 : data_o = 1'b0;
            4928 : data_o = 1'b0;
            4929 : data_o = 1'b0;
            4930 : data_o = 1'b0;
            4931 : data_o = 1'b0;
            4932 : data_o = 1'b0;
            4933 : data_o = 1'b0;
            4934 : data_o = 1'b0;
            4935 : data_o = 1'b0;
            4936 : data_o = 1'b0;
            4937 : data_o = 1'b0;
            4938 : data_o = 1'b0;
            4939 : data_o = 1'b0;
            4940 : data_o = 1'b0;
            4941 : data_o = 1'b0;
            4942 : data_o = 1'b0;
            4943 : data_o = 1'b0;
            4944 : data_o = 1'b0;
            4945 : data_o = 1'b0;
            4946 : data_o = 1'b0;
            4947 : data_o = 1'b0;
            4948 : data_o = 1'b0;
            4949 : data_o = 1'b0;
            4950 : data_o = 1'b0;
            4951 : data_o = 1'b0;
            4952 : data_o = 1'b0;
            4953 : data_o = 1'b1;
            4954 : data_o = 1'b1;
            4955 : data_o = 1'b1;
            4956 : data_o = 1'b1;
            4957 : data_o = 1'b1;
            4958 : data_o = 1'b1;
            4959 : data_o = 1'b1;
            4960 : data_o = 1'b1;
            4961 : data_o = 1'b1;
            4962 : data_o = 1'b1;
            4963 : data_o = 1'b1;
            4964 : data_o = 1'b1;
            4965 : data_o = 1'b1;
            4966 : data_o = 1'b1;
            4967 : data_o = 1'b1;
            4968 : data_o = 1'b1;
            4969 : data_o = 1'b1;
            4970 : data_o = 1'b1;
            4971 : data_o = 1'b1;
            4972 : data_o = 1'b1;
            4973 : data_o = 1'b1;
            4974 : data_o = 1'b1;
            4975 : data_o = 1'b1;
            4976 : data_o = 1'b1;
            4977 : data_o = 1'b1;
            4978 : data_o = 1'b1;
            4979 : data_o = 1'b1;
            4980 : data_o = 1'b1;
            4981 : data_o = 1'b1;
            4982 : data_o = 1'b1;
            4983 : data_o = 1'b1;
            4984 : data_o = 1'b1;
            4985 : data_o = 1'b1;
            4986 : data_o = 1'b1;
            4987 : data_o = 1'b1;
            4988 : data_o = 1'b1;
            4989 : data_o = 1'b1;
            4990 : data_o = 1'b1;
            4991 : data_o = 1'b1;
            4992 : data_o = 1'b1;
            4993 : data_o = 1'b1;
            4994 : data_o = 1'b1;
            4995 : data_o = 1'b1;
            4996 : data_o = 1'b1;
            4997 : data_o = 1'b1;
            4998 : data_o = 1'b1;
            4999 : data_o = 1'b1;
            5000 : data_o = 1'b1;
            5001 : data_o = 1'b1;
            5002 : data_o = 1'b1;
            5003 : data_o = 1'b1;
            5004 : data_o = 1'b1;
            5005 : data_o = 1'b1;
            5006 : data_o = 1'b0;
            5007 : data_o = 1'b0;
            5008 : data_o = 1'b0;
            5009 : data_o = 1'b0;
            5010 : data_o = 1'b0;
            5011 : data_o = 1'b0;
            5012 : data_o = 1'b0;
            5013 : data_o = 1'b0;
            5014 : data_o = 1'b0;
            5015 : data_o = 1'b0;
            5016 : data_o = 1'b0;
            5017 : data_o = 1'b0;
            5018 : data_o = 1'b0;
            5019 : data_o = 1'b0;
            5020 : data_o = 1'b0;
            5021 : data_o = 1'b0;
            5022 : data_o = 1'b0;
            5023 : data_o = 1'b0;
            5024 : data_o = 1'b0;
            5025 : data_o = 1'b0;
            5026 : data_o = 1'b0;
            5027 : data_o = 1'b0;
            5028 : data_o = 1'b0;
            5029 : data_o = 1'b0;
            5030 : data_o = 1'b0;
            5031 : data_o = 1'b0;
            5032 : data_o = 1'b0;
            5033 : data_o = 1'b0;
            5034 : data_o = 1'b0;
            5035 : data_o = 1'b0;
            5036 : data_o = 1'b0;
            5037 : data_o = 1'b0;
            5038 : data_o = 1'b0;
            5039 : data_o = 1'b0;
            5040 : data_o = 1'b0;
            5041 : data_o = 1'b0;
            5042 : data_o = 1'b0;
            5043 : data_o = 1'b0;
            5044 : data_o = 1'b0;
            5045 : data_o = 1'b0;
            5046 : data_o = 1'b0;
            5047 : data_o = 1'b0;
            5048 : data_o = 1'b0;
            5049 : data_o = 1'b0;
            5050 : data_o = 1'b0;
            5051 : data_o = 1'b0;
            5052 : data_o = 1'b0;
            5053 : data_o = 1'b0;
            5054 : data_o = 1'b0;
            5055 : data_o = 1'b0;
            5056 : data_o = 1'b0;
            5057 : data_o = 1'b0;
            5058 : data_o = 1'b0;
            5059 : data_o = 1'b0;
            5060 : data_o = 1'b1;
            5061 : data_o = 1'b1;
            5062 : data_o = 1'b1;
            5063 : data_o = 1'b1;
            5064 : data_o = 1'b1;
            5065 : data_o = 1'b1;
            5066 : data_o = 1'b1;
            5067 : data_o = 1'b1;
            5068 : data_o = 1'b1;
            5069 : data_o = 1'b1;
            5070 : data_o = 1'b1;
            5071 : data_o = 1'b1;
            5072 : data_o = 1'b1;
            5073 : data_o = 1'b1;
            5074 : data_o = 1'b1;
            5075 : data_o = 1'b1;
            5076 : data_o = 1'b1;
            5077 : data_o = 1'b1;
            5078 : data_o = 1'b1;
            5079 : data_o = 1'b1;
            5080 : data_o = 1'b1;
            5081 : data_o = 1'b1;
            5082 : data_o = 1'b1;
            5083 : data_o = 1'b1;
            5084 : data_o = 1'b1;
            5085 : data_o = 1'b1;
            5086 : data_o = 1'b1;
            5087 : data_o = 1'b1;
            5088 : data_o = 1'b1;
            5089 : data_o = 1'b1;
            5090 : data_o = 1'b1;
            5091 : data_o = 1'b1;
            5092 : data_o = 1'b1;
            5093 : data_o = 1'b1;
            5094 : data_o = 1'b1;
            5095 : data_o = 1'b1;
            5096 : data_o = 1'b1;
            5097 : data_o = 1'b1;
            5098 : data_o = 1'b1;
            5099 : data_o = 1'b1;
            5100 : data_o = 1'b1;
            5101 : data_o = 1'b1;
            5102 : data_o = 1'b1;
            5103 : data_o = 1'b1;
            5104 : data_o = 1'b1;
            5105 : data_o = 1'b1;
            5106 : data_o = 1'b1;
            5107 : data_o = 1'b1;
            5108 : data_o = 1'b1;
            5109 : data_o = 1'b1;
            5110 : data_o = 1'b1;
            5111 : data_o = 1'b1;
            5112 : data_o = 1'b1;
            5113 : data_o = 1'b0;
            5114 : data_o = 1'b0;
            5115 : data_o = 1'b0;
            5116 : data_o = 1'b0;
            5117 : data_o = 1'b0;
            5118 : data_o = 1'b0;
            5119 : data_o = 1'b0;
            5120 : data_o = 1'b0;
            5121 : data_o = 1'b0;
            5122 : data_o = 1'b0;
            5123 : data_o = 1'b0;
            5124 : data_o = 1'b0;
            5125 : data_o = 1'b0;
            5126 : data_o = 1'b0;
            5127 : data_o = 1'b0;
            5128 : data_o = 1'b0;
            5129 : data_o = 1'b0;
            5130 : data_o = 1'b0;
            5131 : data_o = 1'b0;
            5132 : data_o = 1'b0;
            5133 : data_o = 1'b0;
            5134 : data_o = 1'b0;
            5135 : data_o = 1'b0;
            5136 : data_o = 1'b0;
            5137 : data_o = 1'b0;
            5138 : data_o = 1'b0;
            5139 : data_o = 1'b0;
            5140 : data_o = 1'b0;
            5141 : data_o = 1'b0;
            5142 : data_o = 1'b0;
            5143 : data_o = 1'b0;
            5144 : data_o = 1'b0;
            5145 : data_o = 1'b0;
            5146 : data_o = 1'b0;
            5147 : data_o = 1'b0;
            5148 : data_o = 1'b0;
            5149 : data_o = 1'b0;
            5150 : data_o = 1'b0;
            5151 : data_o = 1'b0;
            5152 : data_o = 1'b0;
            5153 : data_o = 1'b0;
            5154 : data_o = 1'b0;
            5155 : data_o = 1'b0;
            5156 : data_o = 1'b0;
            5157 : data_o = 1'b0;
            5158 : data_o = 1'b0;
            5159 : data_o = 1'b0;
            5160 : data_o = 1'b0;
            5161 : data_o = 1'b0;
            5162 : data_o = 1'b0;
            5163 : data_o = 1'b0;
            5164 : data_o = 1'b0;
            5165 : data_o = 1'b0;
            5166 : data_o = 1'b0;
            5167 : data_o = 1'b0;
            5168 : data_o = 1'b0;
            5169 : data_o = 1'b1;
            5170 : data_o = 1'b1;
            5171 : data_o = 1'b1;
            5172 : data_o = 1'b1;
            5173 : data_o = 1'b1;
            5174 : data_o = 1'b1;
            5175 : data_o = 1'b1;
            5176 : data_o = 1'b1;
            5177 : data_o = 1'b1;
            5178 : data_o = 1'b1;
            5179 : data_o = 1'b1;
            5180 : data_o = 1'b1;
            5181 : data_o = 1'b1;
            5182 : data_o = 1'b1;
            5183 : data_o = 1'b1;
            5184 : data_o = 1'b1;
            5185 : data_o = 1'b1;
            5186 : data_o = 1'b1;
            5187 : data_o = 1'b1;
            5188 : data_o = 1'b1;
            5189 : data_o = 1'b1;
            5190 : data_o = 1'b1;
            5191 : data_o = 1'b1;
            5192 : data_o = 1'b1;
            5193 : data_o = 1'b1;
            5194 : data_o = 1'b1;
            5195 : data_o = 1'b1;
            5196 : data_o = 1'b1;
            5197 : data_o = 1'b1;
            5198 : data_o = 1'b1;
            5199 : data_o = 1'b1;
            5200 : data_o = 1'b1;
            5201 : data_o = 1'b1;
            5202 : data_o = 1'b1;
            5203 : data_o = 1'b1;
            5204 : data_o = 1'b1;
            5205 : data_o = 1'b1;
            5206 : data_o = 1'b1;
            5207 : data_o = 1'b0;
            5208 : data_o = 1'b0;
            5209 : data_o = 1'b0;
            5210 : data_o = 1'b1;
            5211 : data_o = 1'b1;
            5212 : data_o = 1'b1;
            5213 : data_o = 1'b1;
            5214 : data_o = 1'b1;
            5215 : data_o = 1'b1;
            5216 : data_o = 1'b1;
            5217 : data_o = 1'b1;
            5218 : data_o = 1'b1;
            5219 : data_o = 1'b1;
            5220 : data_o = 1'b0;
            5221 : data_o = 1'b0;
            5222 : data_o = 1'b0;
            5223 : data_o = 1'b0;
            5224 : data_o = 1'b0;
            5225 : data_o = 1'b0;
            5226 : data_o = 1'b0;
            5227 : data_o = 1'b0;
            5228 : data_o = 1'b0;
            5229 : data_o = 1'b0;
            5230 : data_o = 1'b0;
            5231 : data_o = 1'b0;
            5232 : data_o = 1'b0;
            5233 : data_o = 1'b0;
            5234 : data_o = 1'b0;
            5235 : data_o = 1'b0;
            5236 : data_o = 1'b0;
            5237 : data_o = 1'b0;
            5238 : data_o = 1'b0;
            5239 : data_o = 1'b0;
            5240 : data_o = 1'b0;
            5241 : data_o = 1'b0;
            5242 : data_o = 1'b0;
            5243 : data_o = 1'b0;
            5244 : data_o = 1'b0;
            5245 : data_o = 1'b0;
            5246 : data_o = 1'b0;
            5247 : data_o = 1'b0;
            5248 : data_o = 1'b0;
            5249 : data_o = 1'b0;
            5250 : data_o = 1'b0;
            5251 : data_o = 1'b0;
            5252 : data_o = 1'b0;
            5253 : data_o = 1'b0;
            5254 : data_o = 1'b0;
            5255 : data_o = 1'b0;
            5256 : data_o = 1'b0;
            5257 : data_o = 1'b0;
            5258 : data_o = 1'b0;
            5259 : data_o = 1'b0;
            5260 : data_o = 1'b0;
            5261 : data_o = 1'b0;
            5262 : data_o = 1'b0;
            5263 : data_o = 1'b0;
            5264 : data_o = 1'b0;
            5265 : data_o = 1'b0;
            5266 : data_o = 1'b0;
            5267 : data_o = 1'b0;
            5268 : data_o = 1'b0;
            5269 : data_o = 1'b0;
            5270 : data_o = 1'b0;
            5271 : data_o = 1'b0;
            5272 : data_o = 1'b0;
            5273 : data_o = 1'b0;
            5274 : data_o = 1'b0;
            5275 : data_o = 1'b1;
            5276 : data_o = 1'b1;
            5277 : data_o = 1'b1;
            5278 : data_o = 1'b1;
            5279 : data_o = 1'b1;
            5280 : data_o = 1'b1;
            5281 : data_o = 1'b1;
            5282 : data_o = 1'b1;
            5283 : data_o = 1'b1;
            5284 : data_o = 1'b1;
            5285 : data_o = 1'b1;
            5286 : data_o = 1'b1;
            5287 : data_o = 1'b1;
            5288 : data_o = 1'b1;
            5289 : data_o = 1'b1;
            5290 : data_o = 1'b1;
            5291 : data_o = 1'b1;
            5292 : data_o = 1'b1;
            5293 : data_o = 1'b1;
            5294 : data_o = 1'b1;
            5295 : data_o = 1'b1;
            5296 : data_o = 1'b1;
            5297 : data_o = 1'b1;
            5298 : data_o = 1'b1;
            5299 : data_o = 1'b1;
            5300 : data_o = 1'b1;
            5301 : data_o = 1'b1;
            5302 : data_o = 1'b1;
            5303 : data_o = 1'b1;
            5304 : data_o = 1'b1;
            5305 : data_o = 1'b1;
            5306 : data_o = 1'b1;
            5307 : data_o = 1'b1;
            5308 : data_o = 1'b1;
            5309 : data_o = 1'b1;
            5310 : data_o = 1'b1;
            5311 : data_o = 1'b1;
            5312 : data_o = 1'b1;
            5313 : data_o = 1'b1;
            5314 : data_o = 1'b0;
            5315 : data_o = 1'b0;
            5316 : data_o = 1'b0;
            5317 : data_o = 1'b1;
            5318 : data_o = 1'b1;
            5319 : data_o = 1'b1;
            5320 : data_o = 1'b1;
            5321 : data_o = 1'b1;
            5322 : data_o = 1'b1;
            5323 : data_o = 1'b1;
            5324 : data_o = 1'b1;
            5325 : data_o = 1'b0;
            5326 : data_o = 1'b0;
            5327 : data_o = 1'b0;
            5328 : data_o = 1'b0;
            5329 : data_o = 1'b0;
            5330 : data_o = 1'b0;
            5331 : data_o = 1'b0;
            5332 : data_o = 1'b0;
            5333 : data_o = 1'b0;
            5334 : data_o = 1'b0;
            5335 : data_o = 1'b0;
            5336 : data_o = 1'b0;
            5337 : data_o = 1'b0;
            5338 : data_o = 1'b0;
            5339 : data_o = 1'b1;
            5340 : data_o = 1'b1;
            5341 : data_o = 1'b1;
            5342 : data_o = 1'b0;
            5343 : data_o = 1'b0;
            5344 : data_o = 1'b0;
            5345 : data_o = 1'b0;
            5346 : data_o = 1'b0;
            5347 : data_o = 1'b0;
            5348 : data_o = 1'b0;
            5349 : data_o = 1'b0;
            5350 : data_o = 1'b0;
            5351 : data_o = 1'b0;
            5352 : data_o = 1'b0;
            5353 : data_o = 1'b0;
            5354 : data_o = 1'b0;
            5355 : data_o = 1'b0;
            5356 : data_o = 1'b0;
            5357 : data_o = 1'b0;
            5358 : data_o = 1'b0;
            5359 : data_o = 1'b0;
            5360 : data_o = 1'b0;
            5361 : data_o = 1'b0;
            5362 : data_o = 1'b0;
            5363 : data_o = 1'b0;
            5364 : data_o = 1'b0;
            5365 : data_o = 1'b0;
            5366 : data_o = 1'b0;
            5367 : data_o = 1'b0;
            5368 : data_o = 1'b0;
            5369 : data_o = 1'b0;
            5370 : data_o = 1'b0;
            5371 : data_o = 1'b0;
            5372 : data_o = 1'b0;
            5373 : data_o = 1'b0;
            5374 : data_o = 1'b0;
            5375 : data_o = 1'b0;
            5376 : data_o = 1'b0;
            5377 : data_o = 1'b0;
            5378 : data_o = 1'b0;
            5379 : data_o = 1'b0;
            5380 : data_o = 1'b0;
            5381 : data_o = 1'b1;
            5382 : data_o = 1'b1;
            5383 : data_o = 1'b1;
            5384 : data_o = 1'b1;
            5385 : data_o = 1'b1;
            5386 : data_o = 1'b1;
            5387 : data_o = 1'b1;
            5388 : data_o = 1'b1;
            5389 : data_o = 1'b1;
            5390 : data_o = 1'b1;
            5391 : data_o = 1'b1;
            5392 : data_o = 1'b1;
            5393 : data_o = 1'b1;
            5394 : data_o = 1'b1;
            5395 : data_o = 1'b1;
            5396 : data_o = 1'b1;
            5397 : data_o = 1'b1;
            5398 : data_o = 1'b1;
            5399 : data_o = 1'b1;
            5400 : data_o = 1'b1;
            5401 : data_o = 1'b1;
            5402 : data_o = 1'b1;
            5403 : data_o = 1'b1;
            5404 : data_o = 1'b1;
            5405 : data_o = 1'b1;
            5406 : data_o = 1'b1;
            5407 : data_o = 1'b1;
            5408 : data_o = 1'b1;
            5409 : data_o = 1'b1;
            5410 : data_o = 1'b1;
            5411 : data_o = 1'b1;
            5412 : data_o = 1'b1;
            5413 : data_o = 1'b1;
            5414 : data_o = 1'b1;
            5415 : data_o = 1'b1;
            5416 : data_o = 1'b1;
            5417 : data_o = 1'b1;
            5418 : data_o = 1'b0;
            5419 : data_o = 1'b0;
            5420 : data_o = 1'b0;
            5421 : data_o = 1'b0;
            5422 : data_o = 1'b0;
            5423 : data_o = 1'b1;
            5424 : data_o = 1'b1;
            5425 : data_o = 1'b1;
            5426 : data_o = 1'b1;
            5427 : data_o = 1'b1;
            5428 : data_o = 1'b1;
            5429 : data_o = 1'b1;
            5430 : data_o = 1'b1;
            5431 : data_o = 1'b1;
            5432 : data_o = 1'b0;
            5433 : data_o = 1'b0;
            5434 : data_o = 1'b0;
            5435 : data_o = 1'b0;
            5436 : data_o = 1'b0;
            5437 : data_o = 1'b0;
            5438 : data_o = 1'b0;
            5439 : data_o = 1'b0;
            5440 : data_o = 1'b0;
            5441 : data_o = 1'b0;
            5442 : data_o = 1'b0;
            5443 : data_o = 1'b0;
            5444 : data_o = 1'b0;
            5445 : data_o = 1'b0;
            5446 : data_o = 1'b0;
            5447 : data_o = 1'b0;
            5448 : data_o = 1'b0;
            5449 : data_o = 1'b0;
            5450 : data_o = 1'b0;
            5451 : data_o = 1'b0;
            5452 : data_o = 1'b0;
            5453 : data_o = 1'b0;
            5454 : data_o = 1'b0;
            5455 : data_o = 1'b0;
            5456 : data_o = 1'b0;
            5457 : data_o = 1'b0;
            5458 : data_o = 1'b0;
            5459 : data_o = 1'b0;
            5460 : data_o = 1'b0;
            5461 : data_o = 1'b0;
            5462 : data_o = 1'b0;
            5463 : data_o = 1'b0;
            5464 : data_o = 1'b0;
            5465 : data_o = 1'b0;
            5466 : data_o = 1'b0;
            5467 : data_o = 1'b0;
            5468 : data_o = 1'b0;
            5469 : data_o = 1'b0;
            5470 : data_o = 1'b0;
            5471 : data_o = 1'b0;
            5472 : data_o = 1'b0;
            5473 : data_o = 1'b0;
            5474 : data_o = 1'b0;
            5475 : data_o = 1'b0;
            5476 : data_o = 1'b0;
            5477 : data_o = 1'b0;
            5478 : data_o = 1'b0;
            5479 : data_o = 1'b0;
            5480 : data_o = 1'b0;
            5481 : data_o = 1'b0;
            5482 : data_o = 1'b0;
            5483 : data_o = 1'b0;
            5484 : data_o = 1'b0;
            5485 : data_o = 1'b0;
            5486 : data_o = 1'b0;
            5487 : data_o = 1'b1;
            5488 : data_o = 1'b1;
            5489 : data_o = 1'b1;
            5490 : data_o = 1'b1;
            5491 : data_o = 1'b1;
            5492 : data_o = 1'b1;
            5493 : data_o = 1'b1;
            5494 : data_o = 1'b1;
            5495 : data_o = 1'b1;
            5496 : data_o = 1'b1;
            5497 : data_o = 1'b1;
            5498 : data_o = 1'b1;
            5499 : data_o = 1'b1;
            5500 : data_o = 1'b1;
            5501 : data_o = 1'b1;
            5502 : data_o = 1'b1;
            5503 : data_o = 1'b1;
            5504 : data_o = 1'b1;
            5505 : data_o = 1'b1;
            5506 : data_o = 1'b1;
            5507 : data_o = 1'b1;
            5508 : data_o = 1'b1;
            5509 : data_o = 1'b1;
            5510 : data_o = 1'b1;
            5511 : data_o = 1'b1;
            5512 : data_o = 1'b1;
            5513 : data_o = 1'b1;
            5514 : data_o = 1'b1;
            5515 : data_o = 1'b1;
            5516 : data_o = 1'b1;
            5517 : data_o = 1'b1;
            5518 : data_o = 1'b1;
            5519 : data_o = 1'b1;
            5520 : data_o = 1'b1;
            5521 : data_o = 1'b1;
            5522 : data_o = 1'b1;
            5523 : data_o = 1'b1;
            5524 : data_o = 1'b0;
            5525 : data_o = 1'b0;
            5526 : data_o = 1'b0;
            5527 : data_o = 1'b0;
            5528 : data_o = 1'b0;
            5529 : data_o = 1'b1;
            5530 : data_o = 1'b1;
            5531 : data_o = 1'b1;
            5532 : data_o = 1'b1;
            5533 : data_o = 1'b1;
            5534 : data_o = 1'b1;
            5535 : data_o = 1'b1;
            5536 : data_o = 1'b1;
            5537 : data_o = 1'b1;
            5538 : data_o = 1'b1;
            5539 : data_o = 1'b0;
            5540 : data_o = 1'b0;
            5541 : data_o = 1'b0;
            5542 : data_o = 1'b0;
            5543 : data_o = 1'b0;
            5544 : data_o = 1'b0;
            5545 : data_o = 1'b0;
            5546 : data_o = 1'b0;
            5547 : data_o = 1'b0;
            5548 : data_o = 1'b0;
            5549 : data_o = 1'b0;
            5550 : data_o = 1'b0;
            5551 : data_o = 1'b0;
            5552 : data_o = 1'b0;
            5553 : data_o = 1'b0;
            5554 : data_o = 1'b0;
            5555 : data_o = 1'b0;
            5556 : data_o = 1'b0;
            5557 : data_o = 1'b0;
            5558 : data_o = 1'b0;
            5559 : data_o = 1'b0;
            5560 : data_o = 1'b0;
            5561 : data_o = 1'b0;
            5562 : data_o = 1'b0;
            5563 : data_o = 1'b0;
            5564 : data_o = 1'b0;
            5565 : data_o = 1'b0;
            5566 : data_o = 1'b0;
            5567 : data_o = 1'b0;
            5568 : data_o = 1'b0;
            5569 : data_o = 1'b0;
            5570 : data_o = 1'b0;
            5571 : data_o = 1'b0;
            5572 : data_o = 1'b0;
            5573 : data_o = 1'b0;
            5574 : data_o = 1'b0;
            5575 : data_o = 1'b0;
            5576 : data_o = 1'b0;
            5577 : data_o = 1'b0;
            5578 : data_o = 1'b0;
            5579 : data_o = 1'b0;
            5580 : data_o = 1'b0;
            5581 : data_o = 1'b0;
            5582 : data_o = 1'b0;
            5583 : data_o = 1'b0;
            5584 : data_o = 1'b0;
            5585 : data_o = 1'b0;
            5586 : data_o = 1'b0;
            5587 : data_o = 1'b0;
            5588 : data_o = 1'b0;
            5589 : data_o = 1'b0;
            5590 : data_o = 1'b0;
            5591 : data_o = 1'b0;
            5592 : data_o = 1'b0;
            5593 : data_o = 1'b0;
            5594 : data_o = 1'b1;
            5595 : data_o = 1'b1;
            5596 : data_o = 1'b1;
            5597 : data_o = 1'b1;
            5598 : data_o = 1'b1;
            5599 : data_o = 1'b1;
            5600 : data_o = 1'b1;
            5601 : data_o = 1'b1;
            5602 : data_o = 1'b1;
            5603 : data_o = 1'b1;
            5604 : data_o = 1'b1;
            5605 : data_o = 1'b1;
            5606 : data_o = 1'b1;
            5607 : data_o = 1'b1;
            5608 : data_o = 1'b1;
            5609 : data_o = 1'b1;
            5610 : data_o = 1'b1;
            5611 : data_o = 1'b1;
            5612 : data_o = 1'b1;
            5613 : data_o = 1'b1;
            5614 : data_o = 1'b1;
            5615 : data_o = 1'b1;
            5616 : data_o = 1'b1;
            5617 : data_o = 1'b1;
            5618 : data_o = 1'b1;
            5619 : data_o = 1'b1;
            5620 : data_o = 1'b1;
            5621 : data_o = 1'b1;
            5622 : data_o = 1'b1;
            5623 : data_o = 1'b1;
            5624 : data_o = 1'b1;
            5625 : data_o = 1'b1;
            5626 : data_o = 1'b1;
            5627 : data_o = 1'b1;
            5628 : data_o = 1'b1;
            5629 : data_o = 1'b1;
            5630 : data_o = 1'b1;
            5631 : data_o = 1'b1;
            5632 : data_o = 1'b1;
            5633 : data_o = 1'b1;
            5634 : data_o = 1'b1;
            5635 : data_o = 1'b1;
            5636 : data_o = 1'b1;
            5637 : data_o = 1'b1;
            5638 : data_o = 1'b1;
            5639 : data_o = 1'b1;
            5640 : data_o = 1'b1;
            5641 : data_o = 1'b1;
            5642 : data_o = 1'b1;
            5643 : data_o = 1'b1;
            5644 : data_o = 1'b1;
            5645 : data_o = 1'b0;
            5646 : data_o = 1'b0;
            5647 : data_o = 1'b0;
            5648 : data_o = 1'b0;
            5649 : data_o = 1'b0;
            5650 : data_o = 1'b0;
            5651 : data_o = 1'b0;
            5652 : data_o = 1'b0;
            5653 : data_o = 1'b0;
            5654 : data_o = 1'b0;
            5655 : data_o = 1'b0;
            5656 : data_o = 1'b0;
            5657 : data_o = 1'b0;
            5658 : data_o = 1'b0;
            5659 : data_o = 1'b0;
            5660 : data_o = 1'b0;
            5661 : data_o = 1'b0;
            5662 : data_o = 1'b0;
            5663 : data_o = 1'b0;
            5664 : data_o = 1'b0;
            5665 : data_o = 1'b0;
            5666 : data_o = 1'b0;
            5667 : data_o = 1'b0;
            5668 : data_o = 1'b0;
            5669 : data_o = 1'b0;
            5670 : data_o = 1'b0;
            5671 : data_o = 1'b0;
            5672 : data_o = 1'b0;
            5673 : data_o = 1'b0;
            5674 : data_o = 1'b0;
            5675 : data_o = 1'b0;
            5676 : data_o = 1'b0;
            5677 : data_o = 1'b0;
            5678 : data_o = 1'b0;
            5679 : data_o = 1'b0;
            5680 : data_o = 1'b0;
            5681 : data_o = 1'b0;
            5682 : data_o = 1'b0;
            5683 : data_o = 1'b0;
            5684 : data_o = 1'b0;
            5685 : data_o = 1'b0;
            5686 : data_o = 1'b0;
            5687 : data_o = 1'b0;
            5688 : data_o = 1'b0;
            5689 : data_o = 1'b0;
            5690 : data_o = 1'b0;
            5691 : data_o = 1'b0;
            5692 : data_o = 1'b0;
            5693 : data_o = 1'b0;
            5694 : data_o = 1'b0;
            5695 : data_o = 1'b0;
            5696 : data_o = 1'b0;
            5697 : data_o = 1'b0;
            5698 : data_o = 1'b0;
            5699 : data_o = 1'b0;
            5700 : data_o = 1'b0;
            5701 : data_o = 1'b0;
            5702 : data_o = 1'b1;
            5703 : data_o = 1'b1;
            5704 : data_o = 1'b1;
            5705 : data_o = 1'b1;
            5706 : data_o = 1'b1;
            5707 : data_o = 1'b1;
            5708 : data_o = 1'b1;
            5709 : data_o = 1'b1;
            5710 : data_o = 1'b1;
            5711 : data_o = 1'b1;
            5712 : data_o = 1'b1;
            5713 : data_o = 1'b1;
            5714 : data_o = 1'b1;
            5715 : data_o = 1'b1;
            5716 : data_o = 1'b1;
            5717 : data_o = 1'b1;
            5718 : data_o = 1'b1;
            5719 : data_o = 1'b1;
            5720 : data_o = 1'b1;
            5721 : data_o = 1'b1;
            5722 : data_o = 1'b1;
            5723 : data_o = 1'b1;
            5724 : data_o = 1'b1;
            5725 : data_o = 1'b1;
            5726 : data_o = 1'b1;
            5727 : data_o = 1'b1;
            5728 : data_o = 1'b1;
            5729 : data_o = 1'b1;
            5730 : data_o = 1'b1;
            5731 : data_o = 1'b1;
            5732 : data_o = 1'b1;
            5733 : data_o = 1'b1;
            5734 : data_o = 1'b1;
            5735 : data_o = 1'b1;
            5736 : data_o = 1'b1;
            5737 : data_o = 1'b1;
            5738 : data_o = 1'b0;
            5739 : data_o = 1'b0;
            5740 : data_o = 1'b0;
            5741 : data_o = 1'b0;
            5742 : data_o = 1'b0;
            5743 : data_o = 1'b0;
            5744 : data_o = 1'b1;
            5745 : data_o = 1'b1;
            5746 : data_o = 1'b1;
            5747 : data_o = 1'b1;
            5748 : data_o = 1'b1;
            5749 : data_o = 1'b1;
            5750 : data_o = 1'b0;
            5751 : data_o = 1'b0;
            5752 : data_o = 1'b0;
            5753 : data_o = 1'b0;
            5754 : data_o = 1'b0;
            5755 : data_o = 1'b0;
            5756 : data_o = 1'b0;
            5757 : data_o = 1'b0;
            5758 : data_o = 1'b0;
            5759 : data_o = 1'b0;
            5760 : data_o = 1'b0;
            5761 : data_o = 1'b0;
            5762 : data_o = 1'b0;
            5763 : data_o = 1'b0;
            5764 : data_o = 1'b0;
            5765 : data_o = 1'b0;
            5766 : data_o = 1'b0;
            5767 : data_o = 1'b0;
            5768 : data_o = 1'b0;
            5769 : data_o = 1'b0;
            5770 : data_o = 1'b0;
            5771 : data_o = 1'b0;
            5772 : data_o = 1'b0;
            5773 : data_o = 1'b0;
            5774 : data_o = 1'b0;
            5775 : data_o = 1'b0;
            5776 : data_o = 1'b0;
            5777 : data_o = 1'b0;
            5778 : data_o = 1'b0;
            5779 : data_o = 1'b0;
            5780 : data_o = 1'b0;
            5781 : data_o = 1'b0;
            5782 : data_o = 1'b0;
            5783 : data_o = 1'b0;
            5784 : data_o = 1'b0;
            5785 : data_o = 1'b0;
            5786 : data_o = 1'b0;
            5787 : data_o = 1'b0;
            5788 : data_o = 1'b0;
            5789 : data_o = 1'b0;
            5790 : data_o = 1'b0;
            5791 : data_o = 1'b0;
            5792 : data_o = 1'b0;
            5793 : data_o = 1'b0;
            5794 : data_o = 1'b0;
            5795 : data_o = 1'b0;
            5796 : data_o = 1'b0;
            5797 : data_o = 1'b0;
            5798 : data_o = 1'b0;
            5799 : data_o = 1'b0;
            5800 : data_o = 1'b0;
            5801 : data_o = 1'b0;
            5802 : data_o = 1'b0;
            5803 : data_o = 1'b0;
            5804 : data_o = 1'b0;
            5805 : data_o = 1'b0;
            5806 : data_o = 1'b0;
            5807 : data_o = 1'b1;
            5808 : data_o = 1'b1;
            5809 : data_o = 1'b1;
            5810 : data_o = 1'b1;
            5811 : data_o = 1'b1;
            5812 : data_o = 1'b1;
            5813 : data_o = 1'b1;
            5814 : data_o = 1'b1;
            5815 : data_o = 1'b1;
            5816 : data_o = 1'b1;
            5817 : data_o = 1'b1;
            5818 : data_o = 1'b1;
            5819 : data_o = 1'b1;
            5820 : data_o = 1'b1;
            5821 : data_o = 1'b1;
            5822 : data_o = 1'b1;
            5823 : data_o = 1'b1;
            5824 : data_o = 1'b1;
            5825 : data_o = 1'b1;
            5826 : data_o = 1'b1;
            5827 : data_o = 1'b1;
            5828 : data_o = 1'b1;
            5829 : data_o = 1'b1;
            5830 : data_o = 1'b1;
            5831 : data_o = 1'b1;
            5832 : data_o = 1'b1;
            5833 : data_o = 1'b1;
            5834 : data_o = 1'b1;
            5835 : data_o = 1'b1;
            5836 : data_o = 1'b1;
            5837 : data_o = 1'b1;
            5838 : data_o = 1'b1;
            5839 : data_o = 1'b1;
            5840 : data_o = 1'b1;
            5841 : data_o = 1'b1;
            5842 : data_o = 1'b1;
            5843 : data_o = 1'b1;
            5844 : data_o = 1'b1;
            5845 : data_o = 1'b1;
            5846 : data_o = 1'b0;
            5847 : data_o = 1'b0;
            5848 : data_o = 1'b0;
            5849 : data_o = 1'b0;
            5850 : data_o = 1'b0;
            5851 : data_o = 1'b1;
            5852 : data_o = 1'b1;
            5853 : data_o = 1'b1;
            5854 : data_o = 1'b1;
            5855 : data_o = 1'b1;
            5856 : data_o = 1'b1;
            5857 : data_o = 1'b0;
            5858 : data_o = 1'b0;
            5859 : data_o = 1'b0;
            5860 : data_o = 1'b0;
            5861 : data_o = 1'b0;
            5862 : data_o = 1'b0;
            5863 : data_o = 1'b0;
            5864 : data_o = 1'b0;
            5865 : data_o = 1'b0;
            5866 : data_o = 1'b0;
            5867 : data_o = 1'b0;
            5868 : data_o = 1'b0;
            5869 : data_o = 1'b0;
            5870 : data_o = 1'b0;
            5871 : data_o = 1'b0;
            5872 : data_o = 1'b0;
            5873 : data_o = 1'b0;
            5874 : data_o = 1'b0;
            5875 : data_o = 1'b0;
            5876 : data_o = 1'b0;
            5877 : data_o = 1'b0;
            5878 : data_o = 1'b0;
            5879 : data_o = 1'b0;
            5880 : data_o = 1'b0;
            5881 : data_o = 1'b0;
            5882 : data_o = 1'b0;
            5883 : data_o = 1'b0;
            5884 : data_o = 1'b0;
            5885 : data_o = 1'b0;
            5886 : data_o = 1'b0;
            5887 : data_o = 1'b0;
            5888 : data_o = 1'b0;
            5889 : data_o = 1'b0;
            5890 : data_o = 1'b0;
            5891 : data_o = 1'b0;
            5892 : data_o = 1'b0;
            5893 : data_o = 1'b0;
            5894 : data_o = 1'b0;
            5895 : data_o = 1'b0;
            5896 : data_o = 1'b0;
            5897 : data_o = 1'b0;
            5898 : data_o = 1'b0;
            5899 : data_o = 1'b0;
            5900 : data_o = 1'b0;
            5901 : data_o = 1'b0;
            5902 : data_o = 1'b0;
            5903 : data_o = 1'b0;
            5904 : data_o = 1'b0;
            5905 : data_o = 1'b0;
            5906 : data_o = 1'b0;
            5907 : data_o = 1'b0;
            5908 : data_o = 1'b0;
            5909 : data_o = 1'b0;
            5910 : data_o = 1'b0;
            5911 : data_o = 1'b0;
            5912 : data_o = 1'b0;
            5913 : data_o = 1'b0;
            5914 : data_o = 1'b0;
            5915 : data_o = 1'b1;
            5916 : data_o = 1'b1;
            5917 : data_o = 1'b1;
            5918 : data_o = 1'b1;
            5919 : data_o = 1'b1;
            5920 : data_o = 1'b1;
            5921 : data_o = 1'b1;
            5922 : data_o = 1'b1;
            5923 : data_o = 1'b1;
            5924 : data_o = 1'b1;
            5925 : data_o = 1'b1;
            5926 : data_o = 1'b1;
            5927 : data_o = 1'b1;
            5928 : data_o = 1'b1;
            5929 : data_o = 1'b1;
            5930 : data_o = 1'b1;
            5931 : data_o = 1'b1;
            5932 : data_o = 1'b1;
            5933 : data_o = 1'b1;
            5934 : data_o = 1'b1;
            5935 : data_o = 1'b1;
            5936 : data_o = 1'b1;
            5937 : data_o = 1'b1;
            5938 : data_o = 1'b1;
            5939 : data_o = 1'b1;
            5940 : data_o = 1'b1;
            5941 : data_o = 1'b1;
            5942 : data_o = 1'b1;
            5943 : data_o = 1'b1;
            5944 : data_o = 1'b1;
            5945 : data_o = 1'b1;
            5946 : data_o = 1'b1;
            5947 : data_o = 1'b1;
            5948 : data_o = 1'b1;
            5949 : data_o = 1'b1;
            5950 : data_o = 1'b1;
            5951 : data_o = 1'b1;
            5952 : data_o = 1'b1;
            5953 : data_o = 1'b1;
            5954 : data_o = 1'b1;
            5955 : data_o = 1'b1;
            5956 : data_o = 1'b1;
            5957 : data_o = 1'b1;
            5958 : data_o = 1'b1;
            5959 : data_o = 1'b1;
            5960 : data_o = 1'b1;
            5961 : data_o = 1'b1;
            5962 : data_o = 1'b1;
            5963 : data_o = 1'b1;
            5964 : data_o = 1'b1;
            5965 : data_o = 1'b1;
            5966 : data_o = 1'b0;
            5967 : data_o = 1'b0;
            5968 : data_o = 1'b0;
            5969 : data_o = 1'b0;
            5970 : data_o = 1'b0;
            5971 : data_o = 1'b0;
            5972 : data_o = 1'b0;
            5973 : data_o = 1'b0;
            5974 : data_o = 1'b0;
            5975 : data_o = 1'b0;
            5976 : data_o = 1'b0;
            5977 : data_o = 1'b0;
            5978 : data_o = 1'b0;
            5979 : data_o = 1'b0;
            5980 : data_o = 1'b0;
            5981 : data_o = 1'b0;
            5982 : data_o = 1'b0;
            5983 : data_o = 1'b0;
            5984 : data_o = 1'b0;
            5985 : data_o = 1'b0;
            5986 : data_o = 1'b0;
            5987 : data_o = 1'b0;
            5988 : data_o = 1'b0;
            5989 : data_o = 1'b0;
            5990 : data_o = 1'b0;
            5991 : data_o = 1'b0;
            5992 : data_o = 1'b0;
            5993 : data_o = 1'b0;
            5994 : data_o = 1'b0;
            5995 : data_o = 1'b0;
            5996 : data_o = 1'b0;
            5997 : data_o = 1'b0;
            5998 : data_o = 1'b0;
            5999 : data_o = 1'b0;
            6000 : data_o = 1'b0;
            6001 : data_o = 1'b0;
            6002 : data_o = 1'b0;
            6003 : data_o = 1'b0;
            6004 : data_o = 1'b0;
            6005 : data_o = 1'b0;
            6006 : data_o = 1'b0;
            6007 : data_o = 1'b0;
            6008 : data_o = 1'b0;
            6009 : data_o = 1'b0;
            6010 : data_o = 1'b0;
            6011 : data_o = 1'b0;
            6012 : data_o = 1'b0;
            6013 : data_o = 1'b0;
            6014 : data_o = 1'b0;
            6015 : data_o = 1'b0;
            6016 : data_o = 1'b0;
            6017 : data_o = 1'b0;
            6018 : data_o = 1'b0;
            6019 : data_o = 1'b0;
            6020 : data_o = 1'b0;
            6021 : data_o = 1'b0;
            6022 : data_o = 1'b0;
            6023 : data_o = 1'b0;
            6024 : data_o = 1'b1;
            6025 : data_o = 1'b1;
            6026 : data_o = 1'b1;
            6027 : data_o = 1'b1;
            6028 : data_o = 1'b1;
            6029 : data_o = 1'b1;
            6030 : data_o = 1'b1;
            6031 : data_o = 1'b1;
            6032 : data_o = 1'b1;
            6033 : data_o = 1'b1;
            6034 : data_o = 1'b1;
            6035 : data_o = 1'b1;
            6036 : data_o = 1'b1;
            6037 : data_o = 1'b1;
            6038 : data_o = 1'b1;
            6039 : data_o = 1'b1;
            6040 : data_o = 1'b1;
            6041 : data_o = 1'b1;
            6042 : data_o = 1'b1;
            6043 : data_o = 1'b1;
            6044 : data_o = 1'b1;
            6045 : data_o = 1'b1;
            6046 : data_o = 1'b1;
            6047 : data_o = 1'b1;
            6048 : data_o = 1'b1;
            6049 : data_o = 1'b1;
            6050 : data_o = 1'b1;
            6051 : data_o = 1'b1;
            6052 : data_o = 1'b1;
            6053 : data_o = 1'b1;
            6054 : data_o = 1'b1;
            6055 : data_o = 1'b1;
            6056 : data_o = 1'b1;
            6057 : data_o = 1'b1;
            6058 : data_o = 1'b1;
            6059 : data_o = 1'b1;
            6060 : data_o = 1'b1;
            6061 : data_o = 1'b1;
            6062 : data_o = 1'b0;
            6063 : data_o = 1'b0;
            6064 : data_o = 1'b0;
            6065 : data_o = 1'b0;
            6066 : data_o = 1'b0;
            6067 : data_o = 1'b1;
            6068 : data_o = 1'b1;
            6069 : data_o = 1'b1;
            6070 : data_o = 1'b1;
            6071 : data_o = 1'b1;
            6072 : data_o = 1'b0;
            6073 : data_o = 1'b0;
            6074 : data_o = 1'b0;
            6075 : data_o = 1'b0;
            6076 : data_o = 1'b0;
            6077 : data_o = 1'b0;
            6078 : data_o = 1'b0;
            6079 : data_o = 1'b0;
            6080 : data_o = 1'b0;
            6081 : data_o = 1'b0;
            6082 : data_o = 1'b0;
            6083 : data_o = 1'b0;
            6084 : data_o = 1'b0;
            6085 : data_o = 1'b0;
            6086 : data_o = 1'b0;
            6087 : data_o = 1'b0;
            6088 : data_o = 1'b0;
            6089 : data_o = 1'b0;
            6090 : data_o = 1'b0;
            6091 : data_o = 1'b0;
            6092 : data_o = 1'b0;
            6093 : data_o = 1'b0;
            6094 : data_o = 1'b0;
            6095 : data_o = 1'b0;
            6096 : data_o = 1'b0;
            6097 : data_o = 1'b0;
            6098 : data_o = 1'b0;
            6099 : data_o = 1'b0;
            6100 : data_o = 1'b0;
            6101 : data_o = 1'b0;
            6102 : data_o = 1'b0;
            6103 : data_o = 1'b0;
            6104 : data_o = 1'b0;
            6105 : data_o = 1'b0;
            6106 : data_o = 1'b0;
            6107 : data_o = 1'b0;
            6108 : data_o = 1'b0;
            6109 : data_o = 1'b0;
            6110 : data_o = 1'b0;
            6111 : data_o = 1'b0;
            6112 : data_o = 1'b0;
            6113 : data_o = 1'b0;
            6114 : data_o = 1'b0;
            6115 : data_o = 1'b0;
            6116 : data_o = 1'b0;
            6117 : data_o = 1'b0;
            6118 : data_o = 1'b0;
            6119 : data_o = 1'b0;
            6120 : data_o = 1'b0;
            6121 : data_o = 1'b0;
            6122 : data_o = 1'b0;
            6123 : data_o = 1'b0;
            6124 : data_o = 1'b0;
            6125 : data_o = 1'b0;
            6126 : data_o = 1'b0;
            6127 : data_o = 1'b0;
            6128 : data_o = 1'b0;
            6129 : data_o = 1'b0;
            6130 : data_o = 1'b0;
            6131 : data_o = 1'b1;
            6132 : data_o = 1'b1;
            6133 : data_o = 1'b1;
            6134 : data_o = 1'b1;
            6135 : data_o = 1'b1;
            6136 : data_o = 1'b1;
            6137 : data_o = 1'b1;
            6138 : data_o = 1'b1;
            6139 : data_o = 1'b1;
            6140 : data_o = 1'b1;
            6141 : data_o = 1'b1;
            6142 : data_o = 1'b1;
            6143 : data_o = 1'b1;
            6144 : data_o = 1'b1;
            6145 : data_o = 1'b1;
            6146 : data_o = 1'b1;
            6147 : data_o = 1'b1;
            6148 : data_o = 1'b1;
            6149 : data_o = 1'b1;
            6150 : data_o = 1'b1;
            6151 : data_o = 1'b1;
            6152 : data_o = 1'b1;
            6153 : data_o = 1'b1;
            6154 : data_o = 1'b1;
            6155 : data_o = 1'b1;
            6156 : data_o = 1'b1;
            6157 : data_o = 1'b1;
            6158 : data_o = 1'b1;
            6159 : data_o = 1'b1;
            6160 : data_o = 1'b1;
            6161 : data_o = 1'b1;
            6162 : data_o = 1'b1;
            6163 : data_o = 1'b1;
            6164 : data_o = 1'b1;
            6165 : data_o = 1'b1;
            6166 : data_o = 1'b1;
            6167 : data_o = 1'b1;
            6168 : data_o = 1'b1;
            6169 : data_o = 1'b1;
            6170 : data_o = 1'b1;
            6171 : data_o = 1'b1;
            6172 : data_o = 1'b1;
            6173 : data_o = 1'b1;
            6174 : data_o = 1'b1;
            6175 : data_o = 1'b1;
            6176 : data_o = 1'b1;
            6177 : data_o = 1'b1;
            6178 : data_o = 1'b1;
            6179 : data_o = 1'b1;
            6180 : data_o = 1'b1;
            6181 : data_o = 1'b0;
            6182 : data_o = 1'b0;
            6183 : data_o = 1'b0;
            6184 : data_o = 1'b0;
            6185 : data_o = 1'b0;
            6186 : data_o = 1'b0;
            6187 : data_o = 1'b0;
            6188 : data_o = 1'b0;
            6189 : data_o = 1'b0;
            6190 : data_o = 1'b0;
            6191 : data_o = 1'b0;
            6192 : data_o = 1'b0;
            6193 : data_o = 1'b0;
            6194 : data_o = 1'b0;
            6195 : data_o = 1'b0;
            6196 : data_o = 1'b0;
            6197 : data_o = 1'b0;
            6198 : data_o = 1'b0;
            6199 : data_o = 1'b0;
            6200 : data_o = 1'b0;
            6201 : data_o = 1'b0;
            6202 : data_o = 1'b0;
            6203 : data_o = 1'b0;
            6204 : data_o = 1'b0;
            6205 : data_o = 1'b0;
            6206 : data_o = 1'b0;
            6207 : data_o = 1'b0;
            6208 : data_o = 1'b0;
            6209 : data_o = 1'b0;
            6210 : data_o = 1'b0;
            6211 : data_o = 1'b0;
            6212 : data_o = 1'b0;
            6213 : data_o = 1'b0;
            6214 : data_o = 1'b0;
            6215 : data_o = 1'b0;
            6216 : data_o = 1'b0;
            6217 : data_o = 1'b0;
            6218 : data_o = 1'b0;
            6219 : data_o = 1'b0;
            6220 : data_o = 1'b0;
            6221 : data_o = 1'b0;
            6222 : data_o = 1'b0;
            6223 : data_o = 1'b0;
            6224 : data_o = 1'b0;
            6225 : data_o = 1'b0;
            6226 : data_o = 1'b0;
            6227 : data_o = 1'b0;
            6228 : data_o = 1'b0;
            6229 : data_o = 1'b0;
            6230 : data_o = 1'b0;
            6231 : data_o = 1'b0;
            6232 : data_o = 1'b0;
            6233 : data_o = 1'b0;
            6234 : data_o = 1'b0;
            6235 : data_o = 1'b0;
            6236 : data_o = 1'b0;
            6237 : data_o = 1'b0;
            6238 : data_o = 1'b1;
            6239 : data_o = 1'b1;
            6240 : data_o = 1'b1;
            6241 : data_o = 1'b1;
            6242 : data_o = 1'b1;
            6243 : data_o = 1'b1;
            6244 : data_o = 1'b1;
            6245 : data_o = 1'b1;
            6246 : data_o = 1'b1;
            6247 : data_o = 1'b1;
            6248 : data_o = 1'b1;
            6249 : data_o = 1'b1;
            6250 : data_o = 1'b1;
            6251 : data_o = 1'b1;
            6252 : data_o = 1'b1;
            6253 : data_o = 1'b1;
            6254 : data_o = 1'b1;
            6255 : data_o = 1'b1;
            6256 : data_o = 1'b1;
            6257 : data_o = 1'b1;
            6258 : data_o = 1'b1;
            6259 : data_o = 1'b1;
            6260 : data_o = 1'b1;
            6261 : data_o = 1'b1;
            6262 : data_o = 1'b1;
            6263 : data_o = 1'b1;
            6264 : data_o = 1'b1;
            6265 : data_o = 1'b1;
            6266 : data_o = 1'b1;
            6267 : data_o = 1'b1;
            6268 : data_o = 1'b1;
            6269 : data_o = 1'b1;
            6270 : data_o = 1'b1;
            6271 : data_o = 1'b1;
            6272 : data_o = 1'b1;
            6273 : data_o = 1'b1;
            6274 : data_o = 1'b1;
            6275 : data_o = 1'b1;
            6276 : data_o = 1'b1;
            6277 : data_o = 1'b1;
            6278 : data_o = 1'b1;
            6279 : data_o = 1'b1;
            6280 : data_o = 1'b1;
            6281 : data_o = 1'b1;
            6282 : data_o = 1'b1;
            6283 : data_o = 1'b1;
            6284 : data_o = 1'b1;
            6285 : data_o = 1'b1;
            6286 : data_o = 1'b0;
            6287 : data_o = 1'b0;
            6288 : data_o = 1'b0;
            6289 : data_o = 1'b0;
            6290 : data_o = 1'b0;
            6291 : data_o = 1'b0;
            6292 : data_o = 1'b0;
            6293 : data_o = 1'b0;
            6294 : data_o = 1'b0;
            6295 : data_o = 1'b0;
            6296 : data_o = 1'b0;
            6297 : data_o = 1'b0;
            6298 : data_o = 1'b0;
            6299 : data_o = 1'b0;
            6300 : data_o = 1'b0;
            6301 : data_o = 1'b0;
            6302 : data_o = 1'b0;
            6303 : data_o = 1'b0;
            6304 : data_o = 1'b0;
            6305 : data_o = 1'b0;
            6306 : data_o = 1'b0;
            6307 : data_o = 1'b0;
            6308 : data_o = 1'b0;
            6309 : data_o = 1'b0;
            6310 : data_o = 1'b0;
            6311 : data_o = 1'b0;
            6312 : data_o = 1'b0;
            6313 : data_o = 1'b0;
            6314 : data_o = 1'b0;
            6315 : data_o = 1'b0;
            6316 : data_o = 1'b0;
            6317 : data_o = 1'b0;
            6318 : data_o = 1'b0;
            6319 : data_o = 1'b0;
            6320 : data_o = 1'b0;
            6321 : data_o = 1'b0;
            6322 : data_o = 1'b0;
            6323 : data_o = 1'b0;
            6324 : data_o = 1'b0;
            6325 : data_o = 1'b0;
            6326 : data_o = 1'b0;
            6327 : data_o = 1'b0;
            6328 : data_o = 1'b0;
            6329 : data_o = 1'b0;
            6330 : data_o = 1'b0;
            6331 : data_o = 1'b0;
            6332 : data_o = 1'b0;
            6333 : data_o = 1'b0;
            6334 : data_o = 1'b0;
            6335 : data_o = 1'b0;
            6336 : data_o = 1'b0;
            6337 : data_o = 1'b0;
            6338 : data_o = 1'b0;
            6339 : data_o = 1'b0;
            6340 : data_o = 1'b0;
            6341 : data_o = 1'b0;
            6342 : data_o = 1'b0;
            6343 : data_o = 1'b0;
            6344 : data_o = 1'b0;
            6345 : data_o = 1'b0;
            6346 : data_o = 1'b1;
            6347 : data_o = 1'b1;
            6348 : data_o = 1'b1;
            6349 : data_o = 1'b1;
            6350 : data_o = 1'b1;
            6351 : data_o = 1'b1;
            6352 : data_o = 1'b1;
            6353 : data_o = 1'b1;
            6354 : data_o = 1'b1;
            6355 : data_o = 1'b1;
            6356 : data_o = 1'b1;
            6357 : data_o = 1'b1;
            6358 : data_o = 1'b1;
            6359 : data_o = 1'b1;
            6360 : data_o = 1'b1;
            6361 : data_o = 1'b1;
            6362 : data_o = 1'b1;
            6363 : data_o = 1'b1;
            6364 : data_o = 1'b1;
            6365 : data_o = 1'b1;
            6366 : data_o = 1'b1;
            6367 : data_o = 1'b1;
            6368 : data_o = 1'b1;
            6369 : data_o = 1'b1;
            6370 : data_o = 1'b1;
            6371 : data_o = 1'b1;
            6372 : data_o = 1'b1;
            6373 : data_o = 1'b1;
            6374 : data_o = 1'b1;
            6375 : data_o = 1'b1;
            6376 : data_o = 1'b1;
            6377 : data_o = 1'b1;
            6378 : data_o = 1'b1;
            6379 : data_o = 1'b1;
            6380 : data_o = 1'b1;
            6381 : data_o = 1'b1;
            6382 : data_o = 1'b1;
            6383 : data_o = 1'b1;
            6384 : data_o = 1'b1;
            6385 : data_o = 1'b1;
            6386 : data_o = 1'b1;
            6387 : data_o = 1'b1;
            6388 : data_o = 1'b1;
            6389 : data_o = 1'b1;
            6390 : data_o = 1'b1;
            6391 : data_o = 1'b1;
            6392 : data_o = 1'b1;
            6393 : data_o = 1'b0;
            6394 : data_o = 1'b0;
            6395 : data_o = 1'b0;
            6396 : data_o = 1'b0;
            6397 : data_o = 1'b0;
            6398 : data_o = 1'b0;
            6399 : data_o = 1'b0;
            6400 : data_o = 1'b0;
            6401 : data_o = 1'b0;
            6402 : data_o = 1'b0;
            6403 : data_o = 1'b0;
            6404 : data_o = 1'b0;
            6405 : data_o = 1'b0;
            6406 : data_o = 1'b0;
            6407 : data_o = 1'b0;
            6408 : data_o = 1'b0;
            6409 : data_o = 1'b0;
            6410 : data_o = 1'b0;
            6411 : data_o = 1'b0;
            6412 : data_o = 1'b0;
            6413 : data_o = 1'b0;
            6414 : data_o = 1'b0;
            6415 : data_o = 1'b0;
            6416 : data_o = 1'b0;
            6417 : data_o = 1'b0;
            6418 : data_o = 1'b0;
            6419 : data_o = 1'b0;
            6420 : data_o = 1'b0;
            6421 : data_o = 1'b0;
            6422 : data_o = 1'b0;
            6423 : data_o = 1'b0;
            6424 : data_o = 1'b0;
            6425 : data_o = 1'b0;
            6426 : data_o = 1'b0;
            6427 : data_o = 1'b0;
            6428 : data_o = 1'b0;
            6429 : data_o = 1'b0;
            6430 : data_o = 1'b0;
            6431 : data_o = 1'b0;
            6432 : data_o = 1'b0;
            6433 : data_o = 1'b0;
            6434 : data_o = 1'b0;
            6435 : data_o = 1'b0;
            6436 : data_o = 1'b0;
            6437 : data_o = 1'b0;
            6438 : data_o = 1'b0;
            6439 : data_o = 1'b0;
            6440 : data_o = 1'b0;
            6441 : data_o = 1'b0;
            6442 : data_o = 1'b0;
            6443 : data_o = 1'b0;
            6444 : data_o = 1'b0;
            6445 : data_o = 1'b0;
            6446 : data_o = 1'b0;
            6447 : data_o = 1'b0;
            6448 : data_o = 1'b0;
            6449 : data_o = 1'b1;
            6450 : data_o = 1'b1;
            6451 : data_o = 1'b1;
            6452 : data_o = 1'b1;
            6453 : data_o = 1'b1;
            6454 : data_o = 1'b1;
            6455 : data_o = 1'b1;
            6456 : data_o = 1'b1;
            6457 : data_o = 1'b1;
            6458 : data_o = 1'b1;
            6459 : data_o = 1'b1;
            6460 : data_o = 1'b1;
            6461 : data_o = 1'b1;
            6462 : data_o = 1'b1;
            6463 : data_o = 1'b1;
            6464 : data_o = 1'b1;
            6465 : data_o = 1'b1;
            6466 : data_o = 1'b1;
            6467 : data_o = 1'b1;
            6468 : data_o = 1'b1;
            6469 : data_o = 1'b1;
            6470 : data_o = 1'b1;
            6471 : data_o = 1'b1;
            6472 : data_o = 1'b1;
            6473 : data_o = 1'b1;
            6474 : data_o = 1'b1;
            6475 : data_o = 1'b1;
            6476 : data_o = 1'b1;
            6477 : data_o = 1'b1;
            6478 : data_o = 1'b1;
            6479 : data_o = 1'b1;
            6480 : data_o = 1'b1;
            6481 : data_o = 1'b1;
            6482 : data_o = 1'b1;
            6483 : data_o = 1'b1;
            6484 : data_o = 1'b1;
            6485 : data_o = 1'b1;
            6486 : data_o = 1'b1;
            6487 : data_o = 1'b1;
            6488 : data_o = 1'b1;
            6489 : data_o = 1'b1;
            6490 : data_o = 1'b1;
            6491 : data_o = 1'b1;
            6492 : data_o = 1'b1;
            6493 : data_o = 1'b1;
            6494 : data_o = 1'b1;
            6495 : data_o = 1'b1;
            6496 : data_o = 1'b1;
            6497 : data_o = 1'b1;
            6498 : data_o = 1'b1;
            6499 : data_o = 1'b1;
            6500 : data_o = 1'b1;
            6501 : data_o = 1'b1;
            6502 : data_o = 1'b1;
            6503 : data_o = 1'b1;
            6504 : data_o = 1'b1;
            6505 : data_o = 1'b1;
            6506 : data_o = 1'b1;
            6507 : data_o = 1'b1;
            6508 : data_o = 1'b1;
            6509 : data_o = 1'b1;
            6510 : data_o = 1'b1;
            6511 : data_o = 1'b1;
            6512 : data_o = 1'b1;
            6513 : data_o = 1'b1;
            6514 : data_o = 1'b1;
            6515 : data_o = 1'b1;
            6516 : data_o = 1'b1;
            6517 : data_o = 1'b1;
            6518 : data_o = 1'b1;
            6519 : data_o = 1'b1;
            6520 : data_o = 1'b1;
            6521 : data_o = 1'b1;
            6522 : data_o = 1'b1;
            6523 : data_o = 1'b1;
            6524 : data_o = 1'b1;
            6525 : data_o = 1'b1;
            6526 : data_o = 1'b1;
            6527 : data_o = 1'b1;
            6528 : data_o = 1'b1;
            6529 : data_o = 1'b1;
            6530 : data_o = 1'b1;
            6531 : data_o = 1'b1;
            6532 : data_o = 1'b1;
            6533 : data_o = 1'b1;
            6534 : data_o = 1'b1;
            6535 : data_o = 1'b1;
            6536 : data_o = 1'b1;
            6537 : data_o = 1'b1;
            6538 : data_o = 1'b1;
            6539 : data_o = 1'b1;
            6540 : data_o = 1'b1;
            6541 : data_o = 1'b1;
            6542 : data_o = 1'b1;
            6543 : data_o = 1'b1;
            6544 : data_o = 1'b1;
            6545 : data_o = 1'b1;
            6546 : data_o = 1'b1;
            6547 : data_o = 1'b1;
            6548 : data_o = 1'b1;
            6549 : data_o = 1'b1;
            6550 : data_o = 1'b1;
            6551 : data_o = 1'b1;
            6552 : data_o = 1'b1;
            6553 : data_o = 1'b1;
            6554 : data_o = 1'b1;
            6555 : data_o = 1'b1;
            6556 : data_o = 1'b1;
            6557 : data_o = 1'b1;
            6558 : data_o = 1'b1;
            6559 : data_o = 1'b1;
            6560 : data_o = 1'b1;
            6561 : data_o = 1'b1;
            6562 : data_o = 1'b1;
            6563 : data_o = 1'b1;
            6564 : data_o = 1'b1;
            6565 : data_o = 1'b1;
            6566 : data_o = 1'b1;
            6567 : data_o = 1'b1;
            6568 : data_o = 1'b1;
            default: data_o = '0;
        endcase
    end
endmodule
