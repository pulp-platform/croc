module bondpad_70x70 (pad);
	inout pad;
endmodule