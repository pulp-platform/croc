.SUBCKT bondpad_70x70 pad
*.PININFO pad:B
.ENDS
